module calculate (
    input clk,
    input reset,
    input [3:0] key_in,
    output reg [3:0] key_out,
    output reg [4:0] led,
    output reg PointTime,
    output reg [3:0] led_int_Data2,
    output reg [3:0] led_int_Data1,
    output reg [3:0] led_int_Data0
);

    reg [7:0]combvalue;
    reg [3:0]scanvalue;
    reg time1Oms;
    reg [15:0] timecnt;

    always @(posedge time1Oms or negedge reset) //clklow为低频128Hz
    begin
        if(reset == 0)
            begin
                scanvalue <= 1;
                led<=5'b11111;
                combvalue<=0;
            end
        else
            begin
                key_out <= scanvalue;
                case(scanvalue)
                    4'b0001:scanvalue<=4'b0010;
                    4'b0010:scanvalue<=4'b0100;
                    4'b0100:scanvalue<=4'b1000;
                    4'b1000:scanvalue<=4'b0001;
                    default:scanvalue<=4'b0001;
                endcase
                combvalue <={key_in , key_out};
                case(combvalue)
                    8'b00010001 : led <= 5'b11110;//1
                    8'b00100001 : led <= 5'b11101;//2
                    8'b01000001 : led <= 5'b11100;//3
                    8'b00010010 : led <= 5'b11010;//4
                    8'b00100010 : led <= 5'b11001;//5
                    8'b01000010 : led <= 5'b11000;//6
                    8'b00010100 : led <= 5'b10110;//7
                    8'b00100100 : led <= 5'b10101;//8
                    8'b01000100 : led <= 5'b10100;//9
                    8'b00011000 : led <= 5'b10010;//0
                    8'b10000001 : led <= 5'b11011;//X
                    8'b10000010 : led <= 5'b10111;//Y
                    8'b10000100 : led <= 5'b10011;//Z
                    8'b00101000 : led <= 5'b10001;//+
                    8'b01001000 : led <= 5'b10000;//-
                    8'b10001000 : led <= 5'b01111;//=
                    default: led <= 5'b11111;
                endcase
            end
    end


    always @(posedge clk or negedge reset) //clk 为系统时钟信号6MHz
    begin
        if(reset==1'b0) timecnt<=0; //timecnt 为分频计数器， 用来得到lOms 时钟
        else if(timecnt==29999)
            begin
                time1Oms<=~time1Oms; //time1Oms 为lOms 时钟
                timecnt<=0;
            end
        else timecnt<=timecnt+ 1;
    end

    reg [1:0] flag_Cal;
    reg [1:0] flag_Data;
    reg flag_Over;
    reg [3:0] int_Data0;
    reg [3:0] int_Data1;
    reg [6:0] int_Data;
    always @(posedge time1Oms or negedge reset)
    begin
        if(reset == 0)
            begin
                flag_Data <= 0;
                flag_Over <= 0;
                flag_Cal <= 0;
                int_Data0 <= 0;
                int_Data1 <= 0;
                PointTime <= 1;
                led_int_Data2 <= 11;
                int_Data <= 0;
            end
        else 
            begin

                case ({key_in , key_out})
                    8'b00010001://1
                        begin
                            case (flag_Data)
                                0: begin led_int_Data2<=11;int_Data0<=1;int_Data<=1;flag_Data<=1;end
                                2: begin int_Data1<=1;int_Data<=1;flag_Data<=3;end 
                                default: ;
                            endcase
                        end
                    8'b00100001://2
                        begin
                            case (flag_Data)
                                0: begin led_int_Data2<=11;int_Data0<=2;int_Data<=2;flag_Data<=1;end
                                2: begin int_Data1<=2;int_Data<=2;flag_Data<=3;end 
                                default: ;
                            endcase
                        end 
                    8'b01000001://3
                        begin
                            case (flag_Data)
                                0: begin led_int_Data2<=11;int_Data0<=3;int_Data<=3;flag_Data<=1;end
                                2: begin int_Data1<=3;int_Data<=3;flag_Data<=3;end 
                                default: ;
                            endcase
                        end
                    8'b00010010://4
                        begin
                            case (flag_Data)
                                0: begin led_int_Data2<=11;int_Data0<=4;int_Data<=4;flag_Data<=1;end
                                2: begin int_Data1<=4;int_Data<=4;flag_Data<=3;end 
                                default: ;
                            endcase
                        end
                    8'b00100010://5
                        begin
                            case (flag_Data)
                                0: begin led_int_Data2<=11;int_Data0<=5;int_Data<=5;flag_Data<=1;end
                                2: begin int_Data1<=5;int_Data<=5;flag_Data<=3;end 
                                default: ;
                            endcase
                        end
                    8'b01000010://6
                        begin
                            case (flag_Data)
                                0: begin led_int_Data2<=11;int_Data0<=6;int_Data<=6;flag_Data<=1;end
                                2: begin int_Data1<=6;int_Data<=6;flag_Data<=3;end 
                                default: ;
                            endcase
                        end
                    8'b00010100://7
                        begin
                            case (flag_Data)
                                0: begin led_int_Data2<=11;int_Data0<=7;int_Data<=7;flag_Data<=1;end
                                2: begin int_Data1<=7;int_Data<=7;flag_Data<=3;end 
                                default: ;
                            endcase
                        end
                    8'b00100100://8
                        begin
                            case (flag_Data)
                                0: begin led_int_Data2<=11;int_Data0<=8;int_Data<=8;flag_Data<=1;end
                                2: begin int_Data1<=8;int_Data<=8;flag_Data<=3;end 
                                default: ;
                            endcase
                        end
                    8'b01000100://9
                        begin
                            case (flag_Data)
                                0: begin led_int_Data2<=11;int_Data0<=9;int_Data<=9;flag_Data<=1;end
                                2: begin int_Data1<=9;int_Data<=9;flag_Data<=3;end 
                                default: ;
                            endcase
                        end
                    8'b00011000://0
                        begin
                            case (flag_Data)
                                0: begin led_int_Data2<=11;int_Data0<=0;int_Data<=0;flag_Data<=1;end
                                2: begin int_Data1<=0;int_Data<=0;flag_Data<=3;end 
                                default: ;
                            endcase
                        end
                    8'b10000001://X
                        begin
                            if(flag_Data==1) begin
                                flag_Cal <= 3;
                                PointTime <= 0;
                                flag_Data <= 2;
                            end
                        end
                    8'b10000010:;//Y
                    8'b10000100://Z
                        begin
                            flag_Over <= 0;
                            flag_Data <= 0;
                            int_Data0 <= 0;
                            int_Data1 <= 0;
                            PointTime <= 1;
                            led_int_Data2 <= 11;
                            int_Data <= 0;
                        end
                    8'b00101000://+
                        begin
                            if(flag_Data==1) begin
                                flag_Cal <= 1;
                                PointTime <= 1;
                                flag_Data <= 2;
                            end
                        end
                    8'b01001000://-
                        begin
                            if(flag_Data == 1)begin
                                flag_Cal <= 2;
                                PointTime <= 0;
                                flag_Data <= 2;
                            end
                        end
                    8'b10001000://=
                        begin
                            case (flag_Cal)
                                1: begin int_Data<=int_Data0+int_Data1;led_int_Data2<=11;end
                                2: begin
                                    if(int_Data0>=int_Data1)
                                        begin
                                            int_Data<=int_Data0-int_Data1;
                                            led_int_Data2<=11;
                                        end
                                    else
                                        begin
                                            int_Data<=int_Data1-int_Data0;
                                            led_int_Data2 <= 10;
                                        end 
                                end
                                3: begin    
                                case({int_Data0,int_Data1})
                                    8'b0000_0000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0000_0001:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0000_0010:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0000_0011:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0000_0100:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0000_0101:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0000_0110:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0000_0111:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0000_1000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0000_1001:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0001_0000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0001_0001:begin int_Data<=1;led_int_Data2<=11;end
                                    8'b0001_0010:begin int_Data<=2;led_int_Data2<=11;end
                                    8'b0001_0011:begin int_Data<=3;led_int_Data2<=11;end
                                    8'b0001_0100:begin int_Data<=4;led_int_Data2<=11;end
                                    8'b0001_0101:begin int_Data<=5;led_int_Data2<=11;end
                                    8'b0001_0110:begin int_Data<=6;led_int_Data2<=11;end
                                    8'b0001_0111:begin int_Data<=7;led_int_Data2<=11;end
                                    8'b0001_1000:begin int_Data<=8;led_int_Data2<=11;end
                                    8'b0001_1001:begin int_Data<=9;led_int_Data2<=11;end
                                    8'b0010_0000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0010_0001:begin int_Data<=2;led_int_Data2<=11;end
                                    8'b0010_0010:begin int_Data<=4;led_int_Data2<=11;end
                                    8'b0010_0011:begin int_Data<=6;led_int_Data2<=11;end
                                    8'b0010_0100:begin int_Data<=8;led_int_Data2<=11;end
                                    8'b0010_0101:begin int_Data<=10;led_int_Data2<=11;end
                                    8'b0010_0110:begin int_Data<=12;led_int_Data2<=11;end
                                    8'b0010_0111:begin int_Data<=14;led_int_Data2<=11;end
                                    8'b0010_1000:begin int_Data<=16;led_int_Data2<=11;end
                                    8'b0010_1001:begin int_Data<=18;led_int_Data2<=11;end
                                    8'b0011_0000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0011_0001:begin int_Data<=3;led_int_Data2<=11;end
                                    8'b0011_0010:begin int_Data<=6;led_int_Data2<=11;end
                                    8'b0011_0011:begin int_Data<=9;led_int_Data2<=11;end
                                    8'b0011_0100:begin int_Data<=12;led_int_Data2<=11;end
                                    8'b0011_0101:begin int_Data<=15;led_int_Data2<=11;end
                                    8'b0011_0110:begin int_Data<=18;led_int_Data2<=11;end
                                    8'b0011_0111:begin int_Data<=21;led_int_Data2<=11;end
                                    8'b0011_1000:begin int_Data<=24;led_int_Data2<=11;end
                                    8'b0011_1001:begin int_Data<=27;led_int_Data2<=11;end
                                    8'b0100_0000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0100_0001:begin int_Data<=4;led_int_Data2<=11;end
                                    8'b0100_0010:begin int_Data<=8;led_int_Data2<=11;end
                                    8'b0100_0011:begin int_Data<=12;led_int_Data2<=11;end
                                    8'b0100_0100:begin int_Data<=16;led_int_Data2<=11;end
                                    8'b0100_0101:begin int_Data<=20;led_int_Data2<=11;end
                                    8'b0100_0110:begin int_Data<=24;led_int_Data2<=11;end
                                    8'b0100_0111:begin int_Data<=28;led_int_Data2<=11;end
                                    8'b0100_1000:begin int_Data<=32;led_int_Data2<=11;end
                                    8'b0100_1001:begin int_Data<=36;led_int_Data2<=11;end
                                    8'b0101_0000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0101_0001:begin int_Data<=5;led_int_Data2<=11;end
                                    8'b0101_0010:begin int_Data<=10;led_int_Data2<=11;end
                                    8'b0101_0011:begin int_Data<=15;led_int_Data2<=11;end
                                    8'b0101_0100:begin int_Data<=20;led_int_Data2<=11;end
                                    8'b0101_0101:begin int_Data<=25;led_int_Data2<=11;end
                                    8'b0101_0110:begin int_Data<=30;led_int_Data2<=11;end
                                    8'b0101_0111:begin int_Data<=35;led_int_Data2<=11;end
                                    8'b0101_1000:begin int_Data<=40;led_int_Data2<=11;end
                                    8'b0101_1001:begin int_Data<=45;led_int_Data2<=11;end
                                    8'b0110_0000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0110_0001:begin int_Data<=6;led_int_Data2<=11;end
                                    8'b0110_0010:begin int_Data<=12;led_int_Data2<=11;end
                                    8'b0110_0011:begin int_Data<=18;led_int_Data2<=11;end
                                    8'b0110_0100:begin int_Data<=24;led_int_Data2<=11;end
                                    8'b0110_0101:begin int_Data<=30;led_int_Data2<=11;end
                                    8'b0110_0110:begin int_Data<=36;led_int_Data2<=11;end
                                    8'b0110_0111:begin int_Data<=42;led_int_Data2<=11;end
                                    8'b0110_1000:begin int_Data<=48;led_int_Data2<=11;end
                                    8'b0110_1001:begin int_Data<=54;led_int_Data2<=11;end
                                    8'b0111_0000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b0111_0001:begin int_Data<=7;led_int_Data2<=11;end
                                    8'b0111_0010:begin int_Data<=14;led_int_Data2<=11;end
                                    8'b0111_0011:begin int_Data<=21;led_int_Data2<=11;end
                                    8'b0111_0100:begin int_Data<=28;led_int_Data2<=11;end
                                    8'b0111_0101:begin int_Data<=35;led_int_Data2<=11;end
                                    8'b0111_0110:begin int_Data<=42;led_int_Data2<=11;end
                                    8'b0111_0111:begin int_Data<=49;led_int_Data2<=11;end
                                    8'b0111_1000:begin int_Data<=56;led_int_Data2<=11;end
                                    8'b0111_1001:begin int_Data<=63;led_int_Data2<=11;end
                                    8'b1000_0000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b1000_0001:begin int_Data<=8;led_int_Data2<=11;end
                                    8'b1000_0010:begin int_Data<=16;led_int_Data2<=11;end
                                    8'b1000_0011:begin int_Data<=24;led_int_Data2<=11;end
                                    8'b1000_0100:begin int_Data<=32;led_int_Data2<=11;end
                                    8'b1000_0101:begin int_Data<=40;led_int_Data2<=11;end
                                    8'b1000_0110:begin int_Data<=48;led_int_Data2<=11;end
                                    8'b1000_0111:begin int_Data<=56;led_int_Data2<=11;end
                                    8'b1000_1000:begin int_Data<=64;led_int_Data2<=11;end
                                    8'b1000_1001:begin int_Data<=72;led_int_Data2<=11;end
                                    8'b1001_0000:begin int_Data<=0;led_int_Data2<=11;end
                                    8'b1001_0001:begin int_Data<=9;led_int_Data2<=11;end
                                    8'b1001_0010:begin int_Data<=18;led_int_Data2<=11;end
                                    8'b1001_0011:begin int_Data<=27;led_int_Data2<=11;end
                                    8'b1001_0100:begin int_Data<=36;led_int_Data2<=11;end
                                    8'b1001_0101:begin int_Data<=45;led_int_Data2<=11;end
                                    8'b1001_0110:begin int_Data<=54;led_int_Data2<=11;end
                                    8'b1001_0111:begin int_Data<=63;led_int_Data2<=11;end
                                    8'b1001_1000:begin int_Data<=72;led_int_Data2<=11;end
                                    8'b1001_1001:begin int_Data<=81;led_int_Data2<=11;end
                                    endcase
                                end 
                                default: ;
                            endcase
                            PointTime <= 1;
                            flag_Cal <= 0;
                            flag_Data <= 0;
                        end
                    default: ;
                endcase
            end
    end

    always @(time1Oms,reset) begin
        if(reset==0)
            begin
                led_int_Data1<=0;led_int_Data0<=0;
            end
        else
            begin
                if(int_Data >79)begin led_int_Data1<=8;led_int_Data0<=int_Data-80; end
                else if(int_Data > 69) begin led_int_Data1<=7;led_int_Data0<=int_Data-70; end
                else if(int_Data > 59) begin led_int_Data1<=6;led_int_Data0<=int_Data-60; end
                else if(int_Data > 49) begin led_int_Data1<=5;led_int_Data0<=int_Data-50; end
                else if(int_Data > 39) begin led_int_Data1<=4;led_int_Data0<=int_Data-40; end
                else if(int_Data > 29) begin led_int_Data1<=3;led_int_Data0<=int_Data-30; end
                else if(int_Data > 19) begin led_int_Data1<=2;led_int_Data0<=int_Data-20; end
                else if(int_Data > 9) begin led_int_Data1<=1;led_int_Data0<=int_Data-10; end
                else begin led_int_Data1<=0; led_int_Data0 <= int_Data; end
            end
    end

endmodule
