// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri May 13 09:16:57 2022
//
// Verilog Description of module lcd1602
//

module lcd1602 (clk_50m, reset, lcdD, lcdRs, lcdRw, ledEN) /* synthesis syn_module_defined=1 */ ;   // lcd1602.v(1[8:15])
    input clk_50m;   // lcd1602.v(2[11:18])
    input reset;   // lcd1602.v(3[11:16])
    output [7:0]lcdD;   // lcd1602.v(4[18:22])
    output lcdRs;   // lcd1602.v(5[16:21])
    output lcdRw;   // lcd1602.v(6[16:21])
    output ledEN;   // lcd1602.v(7[12:17])
    
    wire clk_50m_c /* synthesis SET_AS_NETWORK=clk_50m_c, is_clock=1 */ ;   // lcd1602.v(2[11:18])
    wire ledEN_c /* synthesis is_clock=1, SET_AS_NETWORK=ledEN_c */ ;   // lcd1602.v(7[12:17])
    
    wire lcdRw_c, n5723, reset_c, lcdRs_c, n6279;
    wire [19:0]cnt;   // lcd1602.v(33[16:19])
    wire [7:0]state;   // lcd1602.v(49[15:20])
    
    wire lcdD_c_7, lcdD_c_6, lcdD_c_5, lcdD_c_4, lcdD_c_3, lcdD_c_2, 
        lcdD_c_1, lcdD_c_0;
    wire [5:0]dispCount;   // lcd1602.v(51[15:24])
    
    wire n5141;
    wire [255:0]dataInBuf;   // lcd1602.v(53[17:26])
    
    wire n6047, n6046, n6044, n5134, n6043, n6041, n5057, n5127, 
        n5120, n6040, n6038, n6037, n6035, n6034, n6032, n6031, 
        n6029, n6028, n3047, n3033, n3040, n5113, n5744, n14, 
        n16, n3649, n6026, n1, n5740, n3006, n3733, n3638, n1_adj_1, 
        n2, ledEN_N_622, n5743;
    wire [5:0]dispCount_5__N_347;
    
    wire lcdRs_N_620, lcdRs_N_619, lcdRs_N_618, n6025, n6276, n6273, 
        n6270, n6267, n6264, n6261, n6258, n6023, n6255, n6252, 
        n6249, n6246, n6243, n6240, n6237, n6234, n6231, n6228, 
        n6225, n6222, n6219, n6216, n6213, n6210, n6207, n6204, 
        n6201, n6198, n6195, n6022, n6192, n6189, n6186, n6183, 
        n6180, n6177, n6174, n6171, n6168, n6165, n6162, n6159, 
        n6156, n6153, n6020, n6150, n6147, n6144, n6141, n6138, 
        n6135, n6132, n6129, n6126, n6123, n6120, n6117, n6114, 
        n6111, n6108, n6105, n6102, n6099, n6096, n6093, n6090, 
        n6087, n6084, n6081, n6078, n6075, n6072, n6069, n6066, 
        n6063, n6060, n6057, n6054, n6051, n6048, n6019, n6045, 
        n6042, n6039, n6036, n6033, n6030, n6027, n6024, n6021, 
        n6018, n6015, n6012, n6009, n6006, n6003, n6000, n5997, 
        n5994, n5991, n5988, n5985, n5982, n5979, n5976, n5973, 
        n5970, n5967, n5964, n4376, n5961, n5958, n5955, n5952, 
        n5949, n5946, n5943, n5940, n5937, n5934, n5931, n5928, 
        n5925, n5922, n5919, n5916, n5913, n5910, n5907, n5904, 
        n5901, n5898, n5895, n5892, n5889, n5886, n5883, n5880, 
        n5877, n5874, n5871, n5868, n5865, n5862, n5859, n5856, 
        n5853, n5850, n5847, n5844, n5841, n5838, n5835, n5832, 
        n5829, n5826, n5823, n5820, n5817, n6017, n5814, n5811, 
        n5808, n5805, n5802, n6016, n5799, n5796, n5793, n5790, 
        n5787, n5784, n5781, n5778, n5106, n5775, n5772, n5769, 
        n5766, n5763, n5760, n5721, n5099, n5757, n5754, n5751, 
        n6014, n5719, n6013, n5748, n36, n5717, n6011, n5745, 
        n6010, n5742, n6008, n6007, n5715, n35, n1_adj_2, n2_adj_3, 
        n100, n101, n102, n103, n104, n105, n2_adj_4, n1_adj_5, 
        lcdRs_N_617, n3117, n34, n14_adj_6, n3000, n5207, n6005, 
        n5209, n6004, n6002, n6001, n5205, n5203, n5999, n32, 
        n5201, n5713, n5199, n5197, n5998, n5224, n5996, n5223, 
        n31, n5222, n5221, n5995, n5218, n5216, n5993, n5214, 
        n5212, n5992, n5990, n5718, n5989, n5987, n5986, n5711, 
        n5258, n5659, n6282, n5210, n5741, lcdRs_N_615, n1845, 
        n5984, n5983, n5981, n30, n29, n5980, n28, n27, n5978, 
        n5977, n26, n5709, n5707, n5737, n5735, n7, n5650, n5975, 
        n5974, n5972, n5971, n5969, n5968, n5966, n5965, n1_adj_7, 
        n2_adj_8, n5963, n5962, n5960, n5092, n24, n5703, n5959, 
        n5957, n5956, n23, n5701, n5954, n5953, n5951, n5950, 
        n5948, n5947, n5945, n5944, n5942, n22, n5699, n21, 
        n5697, n5941, n5939, n5938, n5936, n5085, n5935, n5933, 
        n5932, n5930, n5929, n5927, n5926, n5924, n5923, n5695, 
        n5921, n5920, n5918, n5917, n5693, n5915, n5914, n5912, 
        n4374, n5691, n5911, n5909, n5908, n5906, n5905, n5903, 
        n5902, n5900, n5899, n5897, n5896, n5894, n5893, n5891, 
        n5890, n5888, n5887, n3644, n1_adj_9, n9, n5885, n1_adj_10, 
        n5, n5884, n5882, n5881, n5879, n5878, n5876, n5875, 
        n5873, n6294, n5726, n6293, n1_adj_11, n2_adj_12, n5872, 
        n6291, n5870, n6285, n33, n6290, n5869, n6288, n40, 
        n5867, n6287, n44, n3731, n6286, n5253, n6284, n5250, 
        n5866, n6283, n3753, n6281, n60, n6280, n5248, n3739, 
        n5255, n5246, n5739, n86, n87, n88, n89, n90, n93, 
        n2212, n94, n92, n91, n3637, n2199, n6289, n6292, n3729, 
        n3100, n5864, n2185, n2_adj_13, n3012, n95, n96, n97, 
        n20, n2164, n2163, n2162, n2161, n2160, n2159, n6278, 
        n3054, n98, n99, n9_adj_14, n6277, n6275, n5863, n5727, 
        n6274, n6272, n1_adj_15, n2_adj_16, n9_adj_17, n6271, n5861, 
        n6269, n6268, n6266, n5860, n6265, n6263, n5728, pwr, 
        n5858, n5078, n5725, n6262, n6260, n6259, n6257, n5857, 
        n6256, n6254, n6253, n5855, n5854, n6251, n6250, n1_adj_18, 
        n2_adj_19, n6248, n6247, n5852, n6245, n6244, n5851, n6242, 
        n5849, n6241, n6239, n5848, n5724, n6238, n6236, n5846, 
        n6235, n6233, n6232, n5845, n6230, n6229, n5843, n6227, 
        n6226, n5842, n6224, n6223, n5176, n1_adj_20, n2_adj_21, 
        n1_adj_22, n2_adj_23, n9_adj_24, n1_adj_25, n5840, n5689, 
        n5169, n5071, n5839, n5162, n1_adj_26, n2_adj_27, n9_adj_28, 
        n1_adj_29, n2_adj_30, n6221, n6220, n6218, n6217, n1_adj_31, 
        n2_adj_32, n5837, n1_adj_33, n2_adj_34, n6215, n1_adj_35, 
        n2_adj_36, n9_adj_37, n6214, n5836, n6212, n1_adj_38, n2_adj_39, 
        n9_adj_40, n1_adj_41, n2_adj_42, n6211, n1_adj_43, n2_adj_44, 
        n9_adj_45, n1_adj_46, n2_adj_47, n5687, n1_adj_48, n2_adj_49, 
        n9_adj_50, n5834, n5833, n6209, n6208, n1_adj_51, n2_adj_52, 
        n9_adj_53, n1_adj_54, n2_adj_55, n5831, n6206, n1_adj_56, 
        n2_adj_57, n1_adj_58, n2_adj_59, n9_adj_60, n1_adj_61, n2_adj_62, 
        n9_adj_63, n6205, n5830, n6203, n6202, n1_adj_64, n2_adj_65, 
        n9_adj_66, n1_adj_67, n2_adj_68, n6200, n5828, n5685, n1_adj_69, 
        n2_adj_70, n5827, n1_adj_71, n2_adj_72, n9_adj_73, n1_adj_74, 
        n2_adj_75, n9_adj_76, n6199, n5194, n5825, n1_adj_77, n2_adj_78, 
        n1_adj_79, n2_adj_80, n9_adj_81, n6197, n5824, n1_adj_82, 
        n2_adj_83, n9_adj_84, n1_adj_85, n2_adj_86, n9_adj_87, n1_adj_88, 
        n2_adj_89, n9_adj_90, n1_adj_91, n2_adj_92, n6196, n1_adj_93, 
        n2_adj_94, n5822, n1_adj_95, n2_adj_96, n6194, n1_adj_97, 
        n2_adj_98, n9_adj_99, n6193, n1_adj_100, n2_adj_101, n9_adj_102, 
        n1_adj_103, n2_adj_104, n9_adj_105, n1_adj_106, n2_adj_107, 
        n9_adj_108, n1_adj_109, n2_adj_110, n9_adj_111, n1_adj_112, 
        n2_adj_113, n9_adj_114, n1_adj_115, n2_adj_116, n1_adj_117, 
        n2_adj_118, n9_adj_119, n6191, n6190, n5821, n1_adj_120, 
        n2_adj_121, n9_adj_122, n1_adj_123, n2_adj_124, n9_adj_125, 
        n1_adj_126, n2_adj_127, n9_adj_128, n1_adj_129, n2_adj_130, 
        n9_adj_131, n1_adj_132, n2_adj_133, n9_adj_134, n1_adj_135, 
        n2_adj_136, n1_adj_137, n2_adj_138, n9_adj_139, n5819, n5683, 
        n1_adj_140, n2_adj_141, n9_adj_142, n1_adj_143, n2_adj_144, 
        n9_adj_145, n1_adj_146, n2_adj_147, n9_adj_148, n1_adj_149, 
        n2_adj_150, n9_adj_151, n1_adj_152, n2_adj_153, n9_adj_154, 
        n1_adj_155, n2_adj_156, n6188, n1_adj_157, n2_adj_158, n9_adj_159, 
        n6187, n5818, n6185, n1_adj_160, n2_adj_161, n9_adj_162, 
        n1_adj_163, n2_adj_164, n9_adj_165, n1_adj_166, n2_adj_167, 
        n9_adj_168, n1_adj_169, n2_adj_170, n9_adj_171, n1_adj_172, 
        n2_adj_173, n9_adj_174, n1_adj_175, n2_adj_176, n5816, n1_adj_177, 
        n2_adj_178, n9_adj_179, n6184, n5155, n1_adj_180, n2_adj_181, 
        n9_adj_182, n1_adj_183, n2_adj_184, n9_adj_185, n1_adj_186, 
        n2_adj_187, n9_adj_188, n1_adj_189, n2_adj_190, n9_adj_191, 
        n1_adj_192, n2_adj_193, n9_adj_194, n1_adj_195, n2_adj_196, 
        n6182, n1_adj_197, n2_adj_198, n9_adj_199, n5196, n1_adj_200, 
        n2_adj_201, n9_adj_202, n1_adj_203, n2_adj_204, n9_adj_205, 
        n1_adj_206, n2_adj_207, n9_adj_208, n1_adj_209, n2_adj_210, 
        n9_adj_211, n1_adj_212, n2_adj_213, n9_adj_214, n1_adj_215, 
        n2_adj_216, n1_adj_217, n2_adj_218, n9_adj_219, n5815, n5259, 
        n1_adj_220, n2_adj_221, n9_adj_222, n1_adj_223, n2_adj_224, 
        n9_adj_225, n1_adj_226, n2_adj_227, n9_adj_228, n1_adj_229, 
        n2_adj_230, n9_adj_231, n1_adj_232, n2_adj_233, n9_adj_234, 
        n1_adj_235, n2_adj_236, n1_adj_237, n2_adj_238, n9_adj_239, 
        n6181, n1_adj_240, n2_adj_241, n9_adj_242, n1_adj_243, n2_adj_244, 
        n9_adj_245, n1_adj_246, n2_adj_247, n9_adj_248, n1_adj_249, 
        n2_adj_250, n9_adj_251, n1_adj_252, n2_adj_253, n9_adj_254, 
        n1_adj_255, n2_adj_256, n6179, n1_adj_257, n2_adj_258, n9_adj_259, 
        n5813, n5812, n1_adj_260, n2_adj_261, n5810, n1_adj_262, 
        n2_adj_263, n6178, n1_adj_264, n2_adj_265, n1_adj_266, n2_adj_267, 
        n9_adj_268, n1_adj_269, n2_adj_270, n1_adj_271, n2_adj_272, 
        n6176, n1_adj_273, n2_adj_274, n9_adj_275, n6175, n6173, 
        n5809, n1_adj_276, n2_adj_277, n9_adj_278, n1_adj_279, n2_adj_280, 
        n5807, n1_adj_281, n2_adj_282, n6172, n1_adj_283, n2_adj_284, 
        n9_adj_285, n1_adj_286, n2_adj_287, n1_adj_288, n2_adj_289, 
        n1_adj_290, n2_adj_291, n9_adj_292, n6170, n1_adj_293, n2_adj_294, 
        n6169, n1_adj_295, n2_adj_296, n9_adj_297, n1_adj_298, n2_adj_299, 
        n5806, n1_adj_300, n2_adj_301, n9_adj_302, n1_adj_303, n2_adj_304, 
        n6167, n1_adj_305, n2_adj_306, n1_adj_307, n2_adj_308, n9_adj_309, 
        n5804, n1_adj_310, n2_adj_311, n9_adj_312, n1_adj_313, n2_adj_314, 
        n9_adj_315, n1_adj_316, n2_adj_317, n1_adj_318, n2_adj_319, 
        n9_adj_320, n1_adj_321, n2_adj_322, n6166, n1_adj_323, n2_adj_324, 
        n5803, n1_adj_325, n2_adj_326, n9_adj_327, n6164, n5801, 
        n6163, n1_adj_328, n2_adj_329, n6161, n1_adj_330, n2_adj_331, 
        n1_adj_332, n2_adj_333, n9_adj_334, n1_adj_335, n2_adj_336, 
        n9_adj_337, n1_adj_338, n2_adj_339, n1_adj_340, n2_adj_341, 
        n6160, n1_adj_342, n2_adj_343, n9_adj_344, n6158, n1_adj_345, 
        n2_adj_346, n9_adj_347, n1_adj_348, n2_adj_349, n5800, n1_adj_350, 
        n2_adj_351, n9_adj_352, n1_adj_353, n2_adj_354, n9_adj_355, 
        n1_adj_356, n2_adj_357, n6157, n1_adj_358, n2_adj_359, n1_adj_360, 
        n2_adj_361, n9_adj_362, n6155, n5798, n6154, n1_adj_363, 
        n2_adj_364, n5797, n5257, n6152, n5795, n1_adj_365, n2_adj_366, 
        n6151, n5681, n9_adj_367, n1_adj_368, n2_adj_369, n6149, 
        n5794, n6148, n9_adj_370, n1_adj_371, n2_adj_372, n6146, 
        n5792, n6145, n9_adj_373, n1_adj_374, n2_adj_375, n6143, 
        n5791, n6142, n5789, n1_adj_376, n2_adj_377, n6140, n5788, 
        n6139, n6137, n1_adj_378, n2_adj_379, n5679, n9_adj_380, 
        n6136, n6134, n6133, n6131, n1_adj_381, n2_adj_382, n6130, 
        n5677, n9_adj_383, n1_adj_384, n2_adj_385, n6128, n5786, 
        n6127, n9_adj_386, n1_adj_387, n2_adj_388, n6125, n5785, 
        n6124, n9_adj_389, n1_adj_390, n2_adj_391, n6122, n5783, 
        n6121, n9_adj_392, n1_adj_393, n2_adj_394, n6119, n5782, 
        n6118, n1_adj_395, n2_adj_396, n6116, n5780, n6115, n1_adj_397, 
        n2_adj_398, n5675, n9_adj_399, n6113, n6112, n6110, n5779, 
        n6109, n1_adj_400, n2_adj_401, n6107, n9_adj_402, n6106, 
        n1_adj_403, n2_adj_404, n6104, n5673, n9_adj_405, n1_adj_406, 
        n2_adj_407, n6103, n5777, n6101, n9_adj_408, n1_adj_409, 
        n2_adj_410, n6100, n5776, n6098, n9_adj_411, n1_adj_412, 
        n2_adj_413, n6097, n9_adj_414, n5774, n1_adj_415, n2_adj_416, 
        n6095, n6094, n5773, n1_adj_417, n2_adj_418, n6092, n5671, 
        n9_adj_419, n5148, n6091, n5771, n6089, n5770, n1_adj_420, 
        n2_adj_421, n6088, n5768, n6086, n9_adj_422, n1_adj_423, 
        n2_adj_424, n6085, n5767, n6083, n9_adj_425, n1_adj_426, 
        n2_adj_427, n6082, n5765, n6080, n9_adj_428, n5669, n1_adj_429, 
        n2_adj_430, n6079, n9_adj_431, n5764, n6077, n1_adj_432, 
        n2_adj_433, n6076, n9_adj_434, n5762, n6074, n1_adj_435, 
        n2_adj_436, n6073, n5761, n5759, n6071, n1_adj_437, n2_adj_438, 
        n5667, n9_adj_439, n5064, n5758, n6070, n5665, n1_adj_440, 
        n2_adj_441, n3806, n3805, n9_adj_442, n3804, n1_adj_443, 
        n2_adj_444, n5756, n9_adj_445, n6068, n1_adj_446, n2_adj_447, 
        n5755, n9_adj_448, n1_adj_449, n2_adj_450, n6067, n5753, 
        n9_adj_451, n5752, n1_adj_452, n2_adj_453, n6065, n9_adj_454, 
        n1_adj_455, n2_adj_456, n5750, n6064, n6062, n1_adj_457, 
        n2_adj_458, n5749, n4, n9_adj_459, n5720, n5747, n5734, 
        n4_adj_460, n4_adj_461, n5733, n1_adj_462, n2_adj_463, n5661, 
        n9_adj_464, n6061, n5746, n1_adj_465, n2_adj_466, n6059, 
        n9_adj_467, n6058, n1_adj_468, n2_adj_469, n6056, n9_adj_470, 
        n6055, n5729, n1_adj_471, n2_adj_472, n6053, n9_adj_473, 
        n6052, n1_adj_474, n2_adj_475, n6050, n3800, n9_adj_476, 
        n5230, n1_adj_477, n2_adj_478, n5232, n5235, n1_adj_479, 
        n2_adj_480, n5237, n9_adj_481, n5239, n6049, n5242, n5663, 
        n5244, n1_adj_482;
    
    GND i1 (.X(lcdRw_c));
    OR2 i3196 (.O(n6017), .I0(n6016), .I1(n6015));
    AND2 i3198 (.O(n6019), .I0(lcdRs_N_619), .I1(dataInBuf[157]));
    DFFR lcdRs_53 (.Q(lcdRs_c), .D(lcdRs_N_615), .CLK(ledEN_c), .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR dispCount_i0_i0 (.Q(dispCount[0]), .D(n2159), .CLK(ledEN_c), 
          .CE(n3804), .R(reset_c));   // lcd1602.v(62[14] 139[12])
    OR2 select_163_Select_124_i9 (.O(n9_adj_174), .I0(n2_adj_173), .I1(n1_adj_172));
    OR3 i1_adj_1 (.O(n5681), .I0(n2_adj_324), .I1(n1_adj_323), .I2(state[0]));
    OR2 reduce_nor_181_i1 (.O(n1_adj_482), .I0(state[6]), .I1(state[7]));
    AND2 i2332 (.O(n5155), .I0(n5148), .I1(cnt[15]));
    AND2 select_163_Select_254_i1 (.O(n1_adj_479), .I0(state[7]), .I1(n6275));
    AND2 select_163_Select_124_i2 (.O(n2_adj_173), .I0(state[6]), .I1(dataInBuf[116]));
    OR2 i3118 (.O(n5939), .I0(n5938), .I1(n5937));
    AND2 select_163_Select_253_i1 (.O(n1_adj_477), .I0(state[7]), .I1(n6272));
    OR2 select_163_Select_123_i9 (.O(n9_adj_171), .I0(n2_adj_170), .I1(n1_adj_169));
    AND2 i3120 (.O(n5941), .I0(lcdRs_N_619), .I1(dataInBuf[128]));
    AND2 select_163_Select_252_i1 (.O(n1_adj_474), .I0(state[7]), .I1(n6269));
    AND2 select_163_Select_123_i2 (.O(n2_adj_170), .I0(state[6]), .I1(dataInBuf[115]));
    AND2 select_163_Select_251_i1 (.O(n1_adj_471), .I0(state[7]), .I1(n6266));
    AND2 select_163_Select_250_i1 (.O(n1_adj_468), .I0(state[7]), .I1(n6263));
    AND2 select_163_Select_249_i1 (.O(n1_adj_465), .I0(state[7]), .I1(n6260));
    AND2 select_163_Select_248_i1 (.O(n1_adj_462), .I0(state[7]), .I1(n6257));
    OR2 i3121 (.O(n5942), .I0(n5941), .I1(n5940));
    AND2 i3123 (.O(n5944), .I0(lcdRs_N_619), .I1(dataInBuf[129]));
    AND2 select_163_Select_246_i1 (.O(n1_adj_457), .I0(state[7]), .I1(n6254));
    OR2 select_163_Select_122_i9 (.O(n9_adj_168), .I0(n2_adj_167), .I1(n1_adj_166));
    AND3 i3458 (.O(n6279), .I0(n4376), .I1(n4374), .I2(state[4]));
    DFFR state_FSM_i1 (.Q(state[7]), .D(n5257), .CLK(ledEN_c), .R(reset_c));   // lcd1602.v(63[13] 138[20])
    OBUF lcdD_pad_7 (.O(lcdD[7]), .I0(lcdD_c_7));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    DFF cnt_171__i0 (.Q(cnt[0]), .D(n105), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    AND2 select_163_Select_245_i1 (.O(n1_adj_455), .I0(state[7]), .I1(n6251));
    AND2 select_163_Select_122_i2 (.O(n2_adj_167), .I0(state[6]), .I1(dataInBuf[114]));
    AND2 select_163_Select_244_i1 (.O(n1_adj_452), .I0(state[7]), .I1(n6248));
    OR2 select_163_Select_121_i9 (.O(n9_adj_165), .I0(n2_adj_164), .I1(n1_adj_163));
    AND2 select_163_Select_243_i1 (.O(n1_adj_449), .I0(state[7]), .I1(n6245));
    AND2 select_163_Select_242_i1 (.O(n1_adj_446), .I0(state[7]), .I1(n6242));
    OR2 select_163_Select_217_i9 (.O(n9_adj_386), .I0(n2_adj_385), .I1(n1_adj_384));
    AND2 select_163_Select_121_i2 (.O(n2_adj_164), .I0(state[6]), .I1(dataInBuf[113]));
    OR2 select_163_Select_120_i9 (.O(n9_adj_162), .I0(n2_adj_161), .I1(n1_adj_160));
    AND2 select_163_Select_120_i2 (.O(n2_adj_161), .I0(state[6]), .I1(dataInBuf[112]));
    AND2 select_163_Select_241_i1 (.O(n1_adj_443), .I0(state[7]), .I1(n6239));
    OR2 i3124 (.O(n5945), .I0(n5944), .I1(n5943));
    AND2 select_163_Select_240_i1 (.O(n1_adj_440), .I0(state[7]), .I1(n6236));
    AND2 select_163_Select_238_i1 (.O(n1_adj_437), .I0(state[7]), .I1(n6233));
    OR2 select_163_Select_216_i9 (.O(n9_adj_383), .I0(n2_adj_382), .I1(n1_adj_381));
    AND2 select_163_Select_237_i1 (.O(n1_adj_435), .I0(state[7]), .I1(n6230));
    AND2 i1555 (.O(n2164), .I0(n2185), .I1(dispCount_5__N_347[5]));
    AND2 i3417 (.O(n6238), .I0(lcdRs_N_619), .I1(dataInBuf[241]));
    AND2 select_163_Select_236_i1 (.O(n1_adj_432), .I0(state[7]), .I1(n6227));
    OR2 select_163_Select_118_i9 (.O(n9_adj_159), .I0(n2_adj_158), .I1(n1_adj_157));
    AND2 select_163_Select_235_i1 (.O(n1_adj_429), .I0(state[7]), .I1(n6224));
    AND2 select_163_Select_234_i1 (.O(n1_adj_426), .I0(state[7]), .I1(n6221));
    AND2 select_163_Select_118_i2 (.O(n2_adj_158), .I0(state[6]), .I1(dataInBuf[110]));
    AND2 select_163_Select_117_i2 (.O(n2_adj_156), .I0(state[6]), .I1(dataInBuf[109]));
    AND2 select_163_Select_233_i1 (.O(n1_adj_423), .I0(state[7]), .I1(n6218));
    OR2 select_163_Select_116_i9 (.O(n9_adj_154), .I0(n2_adj_153), .I1(n1_adj_152));
    AND2 select_163_Select_232_i1 (.O(n1_adj_420), .I0(state[7]), .I1(n6215));
    AND2 select_163_Select_116_i2 (.O(n2_adj_153), .I0(state[6]), .I1(dataInBuf[108]));
    OR2 select_163_Select_115_i9 (.O(n9_adj_151), .I0(n2_adj_150), .I1(n1_adj_149));
    AND2 select_163_Select_230_i1 (.O(n1_adj_417), .I0(state[7]), .I1(n6212));
    AND2 select_163_Select_115_i2 (.O(n2_adj_150), .I0(state[6]), .I1(dataInBuf[107]));
    OR2 select_163_Select_114_i9 (.O(n9_adj_148), .I0(n2_adj_147), .I1(n1_adj_146));
    AND2 select_163_Select_114_i2 (.O(n2_adj_147), .I0(state[6]), .I1(dataInBuf[106]));
    AND2 select_163_Select_229_i1 (.O(n1_adj_415), .I0(state[7]), .I1(n6209));
    AND2 select_163_Select_228_i1 (.O(n1_adj_412), .I0(state[7]), .I1(n6206));
    AND2 select_163_Select_227_i1 (.O(n1_adj_409), .I0(state[7]), .I1(n6203));
    OR2 select_163_Select_113_i9 (.O(n9_adj_145), .I0(n2_adj_144), .I1(n1_adj_143));
    AND2 select_163_Select_113_i2 (.O(n2_adj_144), .I0(state[6]), .I1(dataInBuf[105]));
    OR2 select_163_Select_112_i9 (.O(n9_adj_142), .I0(n2_adj_141), .I1(n1_adj_140));
    AND2 select_163_Select_226_i1 (.O(n1_adj_406), .I0(state[7]), .I1(n6200));
    AND2 select_163_Select_225_i1 (.O(n1_adj_403), .I0(state[7]), .I1(n6197));
    AND2 select_163_Select_112_i2 (.O(n2_adj_141), .I0(state[6]), .I1(dataInBuf[104]));
    AND2 select_163_Select_224_i1 (.O(n1_adj_400), .I0(state[7]), .I1(n6194));
    OR2 select_163_Select_110_i9 (.O(n9_adj_139), .I0(n2_adj_138), .I1(n1_adj_137));
    AND2 select_163_Select_222_i1 (.O(n1_adj_397), .I0(state[7]), .I1(n6191));
    AND2 select_163_Select_110_i2 (.O(n2_adj_138), .I0(state[6]), .I1(dataInBuf[102]));
    AND2 i3126 (.O(n5947), .I0(lcdRs_N_619), .I1(dataInBuf[130]));
    AND2 select_163_Select_221_i1 (.O(n1_adj_395), .I0(state[7]), .I1(n6188));
    AND2 select_163_Select_220_i1 (.O(n1_adj_393), .I0(state[7]), .I1(n6185));
    OR3 i2 (.O(n5250), .I0(n1_adj_56), .I1(state[0]), .I2(n2_adj_57));
    AND2 select_163_Select_219_i1 (.O(n1_adj_390), .I0(state[7]), .I1(n6182));
    AND2 select_163_Select_218_i1 (.O(n1_adj_387), .I0(state[7]), .I1(n6179));
    AND2 select_163_Select_109_i2 (.O(n2_adj_136), .I0(state[6]), .I1(dataInBuf[101]));
    OR2 select_163_Select_108_i9 (.O(n9_adj_134), .I0(n2_adj_133), .I1(n1_adj_132));
    AND2 select_163_Select_108_i2 (.O(n2_adj_133), .I0(state[6]), .I1(dataInBuf[100]));
    OR2 select_163_Select_107_i9 (.O(n9_adj_131), .I0(n2_adj_130), .I1(n1_adj_129));
    AND2 select_163_Select_217_i1 (.O(n1_adj_384), .I0(state[7]), .I1(n6176));
    AND2 select_163_Select_216_i1 (.O(n1_adj_381), .I0(state[7]), .I1(n6173));
    AND2 select_163_Select_107_i2 (.O(n2_adj_130), .I0(state[6]), .I1(dataInBuf[99]));
    OR2 select_163_Select_106_i9 (.O(n9_adj_128), .I0(n2_adj_127), .I1(n1_adj_126));
    AND2 select_163_Select_214_i1 (.O(n1_adj_378), .I0(state[7]), .I1(n6170));
    AND2 select_163_Select_106_i2 (.O(n2_adj_127), .I0(state[6]), .I1(dataInBuf[98]));
    AND2 select_163_Select_213_i1 (.O(n1_adj_376), .I0(state[7]), .I1(n6167));
    AND2 select_163_Select_212_i1 (.O(n1_adj_374), .I0(state[7]), .I1(n6164));
    OR2 select_163_Select_105_i9 (.O(n9_adj_125), .I0(n2_adj_124), .I1(n1_adj_123));
    AND2 select_163_Select_105_i2 (.O(n2_adj_124), .I0(state[6]), .I1(dataInBuf[97]));
    AND2 select_163_Select_211_i1 (.O(n1_adj_371), .I0(state[7]), .I1(n6161));
    AND2 select_163_Select_210_i1 (.O(n1_adj_368), .I0(state[7]), .I1(n6158));
    OR2 select_163_Select_104_i9 (.O(n9_adj_122), .I0(n2_adj_121), .I1(n1_adj_120));
    AND2 select_163_Select_104_i2 (.O(n2_adj_121), .I0(state[6]), .I1(dataInBuf[96]));
    AND2 select_163_Select_209_i1 (.O(n1_adj_365), .I0(state[7]), .I1(n6155));
    AND2 select_163_Select_208_i1 (.O(n1_adj_363), .I0(state[7]), .I1(n6152));
    AND2 select_163_Select_206_i1 (.O(n1_adj_360), .I0(state[7]), .I1(n6149));
    OR2 i3127 (.O(n5948), .I0(n5947), .I1(n5946));
    OR2 select_163_Select_102_i9 (.O(n9_adj_119), .I0(n2_adj_118), .I1(n1_adj_117));
    AND2 select_163_Select_205_i1 (.O(n1_adj_358), .I0(state[7]), .I1(n6146));
    AND2 select_163_Select_102_i2 (.O(n2_adj_118), .I0(state[6]), .I1(dataInBuf[94]));
    AND2 select_163_Select_101_i2 (.O(n2_adj_116), .I0(state[6]), .I1(dataInBuf[93]));
    OR2 select_163_Select_100_i9 (.O(n9_adj_114), .I0(n2_adj_113), .I1(n1_adj_112));
    AND2 select_163_Select_204_i1 (.O(n1_adj_356), .I0(state[7]), .I1(n6143));
    AND2 select_163_Select_203_i1 (.O(n1_adj_353), .I0(state[7]), .I1(n6140));
    AND2 select_163_Select_202_i1 (.O(n1_adj_350), .I0(state[7]), .I1(n6137));
    AND2 select_163_Select_201_i1 (.O(n1_adj_348), .I0(state[7]), .I1(n6134));
    AND2 select_163_Select_200_i1 (.O(n1_adj_345), .I0(state[7]), .I1(n6131));
    AND2 select_163_Select_100_i2 (.O(n2_adj_113), .I0(state[6]), .I1(dataInBuf[92]));
    OR2 select_163_Select_99_i9 (.O(n9_adj_111), .I0(n2_adj_110), .I1(n1_adj_109));
    AND2 select_163_Select_198_i1 (.O(n1_adj_342), .I0(state[7]), .I1(n6128));
    AND2 select_163_Select_197_i1 (.O(n1_adj_340), .I0(state[7]), .I1(n6125));
    AND2 select_163_Select_99_i2 (.O(n2_adj_110), .I0(state[6]), .I1(dataInBuf[91]));
    OR2 select_163_Select_98_i9 (.O(n9_adj_108), .I0(n2_adj_107), .I1(n1_adj_106));
    AND2 select_163_Select_196_i1 (.O(n1_adj_338), .I0(state[7]), .I1(n6122));
    AND2 select_163_Select_98_i2 (.O(n2_adj_107), .I0(state[6]), .I1(dataInBuf[90]));
    AND2 select_163_Select_195_i1 (.O(n1_adj_335), .I0(state[7]), .I1(n6119));
    OR2 select_163_Select_97_i9 (.O(n9_adj_105), .I0(n2_adj_104), .I1(n1_adj_103));
    AND2 select_163_Select_194_i1 (.O(n1_adj_332), .I0(state[7]), .I1(n6116));
    AND2 select_163_Select_97_i2 (.O(n2_adj_104), .I0(state[6]), .I1(dataInBuf[89]));
    OR2 select_163_Select_96_i9 (.O(n9_adj_102), .I0(n2_adj_101), .I1(n1_adj_100));
    AND2 select_163_Select_193_i1 (.O(n1_adj_330), .I0(state[7]), .I1(n6113));
    AND2 select_163_Select_192_i1 (.O(n1_adj_328), .I0(state[7]), .I1(n6110));
    INV i2916 (.O(n5737), .I0(n3644));
    AND2 select_163_Select_96_i2 (.O(n2_adj_101), .I0(state[6]), .I1(dataInBuf[88]));
    AND2 i3129 (.O(n5950), .I0(lcdRs_N_619), .I1(dataInBuf[131]));
    DFF clkhz_52 (.Q(ledEN_c), .D(ledEN_N_622), .CLK(clk_50m_c));   // lcd1602.v(35[12] 45[8])
    OR2 select_163_Select_94_i9 (.O(n9_adj_99), .I0(n2_adj_98), .I1(n1_adj_97));
    OR2 i3199 (.O(n6020), .I0(n6019), .I1(n6018));
    AND2 select_163_Select_190_i1 (.O(n1_adj_325), .I0(state[7]), .I1(n6107));
    AND2 select_163_Select_94_i2 (.O(n2_adj_98), .I0(state[6]), .I1(dataInBuf[86]));
    AND2 select_163_Select_93_i2 (.O(n2_adj_96), .I0(state[6]), .I1(dataInBuf[85]));
    AND2 select_163_Select_189_i1 (.O(n1_adj_323), .I0(state[7]), .I1(n6104));
    AND2 select_163_Select_188_i1 (.O(n1_adj_321), .I0(state[7]), .I1(n6101));
    AND2 select_163_Select_216_i2 (.O(n2_adj_382), .I0(state[6]), .I1(dataInBuf[208]));
    OR2 i3130 (.O(n5951), .I0(n5950), .I1(n5949));
    AND2 select_163_Select_92_i2 (.O(n2_adj_94), .I0(state[6]), .I1(dataInBuf[84]));
    OR3 i2_adj_2 (.O(n5221), .I0(n1_adj_279), .I1(n2_adj_280), .I2(state[0]));
    AND2 select_163_Select_187_i1 (.O(n1_adj_318), .I0(state[7]), .I1(n6098));
    AND2 select_163_Select_186_i1 (.O(n1_adj_316), .I0(state[7]), .I1(n6095));
    AND2 select_163_Select_185_i1 (.O(n1_adj_313), .I0(state[7]), .I1(n6092));
    IBUF reset_pad (.O(reset_c), .I0(reset));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(186[8:12])
    AND2 select_163_Select_91_i2 (.O(n2_adj_92), .I0(state[6]), .I1(dataInBuf[83]));
    OR2 select_163_Select_90_i9 (.O(n9_adj_90), .I0(n2_adj_89), .I1(n1_adj_88));
    AND2 select_163_Select_90_i2 (.O(n2_adj_89), .I0(state[6]), .I1(dataInBuf[82]));
    AND2 select_163_Select_184_i1 (.O(n1_adj_310), .I0(state[7]), .I1(n6089));
    OR2 select_163_Select_89_i9 (.O(n9_adj_87), .I0(n2_adj_86), .I1(n1_adj_85));
    AND2 select_163_Select_182_i1 (.O(n1_adj_307), .I0(state[7]), .I1(n6086));
    DFF cnt_171__i19 (.Q(cnt[19]), .D(n86), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    AND2 select_163_Select_89_i2 (.O(n2_adj_86), .I0(state[6]), .I1(dataInBuf[81]));
    OR2 select_163_Select_88_i9 (.O(n9_adj_84), .I0(n2_adj_83), .I1(n1_adj_82));
    AND2 select_163_Select_88_i2 (.O(n2_adj_83), .I0(state[6]), .I1(dataInBuf[80]));
    AND2 select_163_Select_181_i1 (.O(n1_adj_305), .I0(state[7]), .I1(n6083));
    AND2 select_163_Select_180_i1 (.O(n1_adj_303), .I0(state[7]), .I1(n6080));
    AND2 select_163_Select_179_i1 (.O(n1_adj_300), .I0(state[7]), .I1(n6077));
    OR2 select_163_Select_86_i9 (.O(n9_adj_81), .I0(n2_adj_80), .I1(n1_adj_79));
    AND2 select_163_Select_178_i1 (.O(n1_adj_298), .I0(state[7]), .I1(n6074));
    AND2 select_163_Select_177_i1 (.O(n1_adj_295), .I0(state[7]), .I1(n6071));
    AND2 select_163_Select_176_i1 (.O(n1_adj_293), .I0(state[7]), .I1(n6068));
    AND2 select_163_Select_86_i2 (.O(n2_adj_80), .I0(state[6]), .I1(dataInBuf[78]));
    AND2 i3132 (.O(n5953), .I0(lcdRs_N_619), .I1(dataInBuf[132]));
    AND2 select_163_Select_85_i2 (.O(n2_adj_78), .I0(state[6]), .I1(dataInBuf[77]));
    OR2 i3133 (.O(n5954), .I0(n5953), .I1(n5952));
    OR2 select_163_Select_82_i9 (.O(n9_adj_76), .I0(n2_adj_75), .I1(n1_adj_74));
    AND2 select_163_Select_174_i1 (.O(n1_adj_290), .I0(state[7]), .I1(n6065));
    AND2 select_163_Select_173_i1 (.O(n1_adj_288), .I0(state[7]), .I1(n6062));
    AND2 select_163_Select_82_i2 (.O(n2_adj_75), .I0(state[6]), .I1(dataInBuf[74]));
    AND2 select_163_Select_172_i1 (.O(n1_adj_286), .I0(state[7]), .I1(n6059));
    OR2 i3292 (.O(n6113), .I0(n6112), .I1(n6111));
    AND2 select_163_Select_171_i1 (.O(n1_adj_283), .I0(state[7]), .I1(n6056));
    OR2 select_163_Select_81_i9 (.O(n9_adj_73), .I0(n2_adj_72), .I1(n1_adj_71));
    AND2 select_163_Select_81_i2 (.O(n2_adj_72), .I0(state[6]), .I1(dataInBuf[73]));
    AND2 select_163_Select_170_i1 (.O(n1_adj_281), .I0(state[7]), .I1(n6053));
    OR3 i2_adj_3 (.O(n5253), .I0(n1_adj_29), .I1(state[0]), .I2(n2_adj_30));
    AND2 select_163_Select_169_i1 (.O(n1_adj_279), .I0(state[7]), .I1(n6050));
    AND2 select_163_Select_80_i2 (.O(n2_adj_70), .I0(state[6]), .I1(dataInBuf[72]));
    AND2 i3135 (.O(n5956), .I0(lcdRs_N_619), .I1(dataInBuf[133]));
    AND2 select_163_Select_168_i1 (.O(n1_adj_276), .I0(state[7]), .I1(n6047));
    AND2 i3201 (.O(n6022), .I0(lcdRs_N_619), .I1(dataInBuf[158]));
    AND2 select_163_Select_166_i1 (.O(n1_adj_273), .I0(state[7]), .I1(n6044));
    AND2 i2283 (.O(n5106), .I0(n5099), .I1(cnt[8]));
    AND2 select_163_Select_78_i2 (.O(n2_adj_68), .I0(state[6]), .I1(dataInBuf[70]));
    AND2 select_163_Select_165_i1 (.O(n1_adj_271), .I0(state[7]), .I1(n6041));
    AND2 select_163_Select_164_i1 (.O(n1_adj_269), .I0(state[7]), .I1(n6038));
    OR2 select_163_Select_77_i9 (.O(n9_adj_66), .I0(n2_adj_65), .I1(n1_adj_64));
    AND2 select_163_Select_77_i2 (.O(n2_adj_65), .I0(state[6]), .I1(dataInBuf[69]));
    AND2 select_163_Select_163_i1 (.O(n1_adj_266), .I0(state[7]), .I1(n6035));
    AND2 select_163_Select_162_i1 (.O(n1_adj_264), .I0(state[7]), .I1(n6032));
    AND2 select_163_Select_161_i1 (.O(n1_adj_262), .I0(state[7]), .I1(n6029));
    AND2 select_163_Select_160_i1 (.O(n1_adj_260), .I0(state[7]), .I1(n6026));
    OR2 select_163_Select_74_i9 (.O(n9_adj_63), .I0(n2_adj_62), .I1(n1_adj_61));
    AND2 select_163_Select_74_i2 (.O(n2_adj_62), .I0(state[6]), .I1(dataInBuf[66]));
    AND2 select_163_Select_158_i1 (.O(n1_adj_257), .I0(state[7]), .I1(n6023));
    AND2 select_163_Select_157_i1 (.O(n1_adj_255), .I0(state[7]), .I1(n6020));
    OR2 select_163_Select_73_i9 (.O(n9_adj_60), .I0(n2_adj_59), .I1(n1_adj_58));
    AND2 select_163_Select_73_i2 (.O(n2_adj_59), .I0(state[6]), .I1(dataInBuf[65]));
    AND2 select_163_Select_156_i1 (.O(n1_adj_252), .I0(state[7]), .I1(n6017));
    OR2 i3136 (.O(n5957), .I0(n5956), .I1(n5955));
    AND2 select_163_Select_155_i1 (.O(n1_adj_249), .I0(state[7]), .I1(n6014));
    AND2 select_163_Select_154_i1 (.O(n1_adj_246), .I0(state[7]), .I1(n6011));
    AND2 select_163_Select_153_i1 (.O(n1_adj_243), .I0(state[7]), .I1(n6008));
    OR2 i1_adj_4 (.O(n4), .I0(state[0]), .I1(n5723));
    AND2 select_163_Select_72_i2 (.O(n2_adj_57), .I0(state[6]), .I1(dataInBuf[64]));
    AND2 select_163_Select_152_i1 (.O(n1_adj_240), .I0(state[7]), .I1(n6005));
    AND2 select_163_Select_150_i1 (.O(n1_adj_237), .I0(state[7]), .I1(n6002));
    AND2 select_163_Select_70_i2 (.O(n2_adj_55), .I0(state[6]), .I1(dataInBuf[62]));
    OR2 select_163_Select_69_i9 (.O(n9_adj_53), .I0(n2_adj_52), .I1(n1_adj_51));
    AND2 select_163_Select_69_i2 (.O(n2_adj_52), .I0(state[6]), .I1(dataInBuf[61]));
    AND2 select_163_Select_149_i1 (.O(n1_adj_235), .I0(state[7]), .I1(n5999));
    AND2 select_163_Select_148_i1 (.O(n1_adj_232), .I0(state[7]), .I1(n5996));
    AND2 i3138 (.O(n5959), .I0(lcdRs_N_619), .I1(dataInBuf[134]));
    OR2 select_163_Select_66_i9 (.O(n9_adj_50), .I0(n2_adj_49), .I1(n1_adj_48));
    AND2 select_163_Select_147_i1 (.O(n1_adj_229), .I0(state[7]), .I1(n5993));
    AND2 select_163_Select_146_i1 (.O(n1_adj_226), .I0(state[7]), .I1(n5990));
    AND2 select_163_Select_145_i1 (.O(n1_adj_223), .I0(state[7]), .I1(n5987));
    AND2 select_163_Select_144_i1 (.O(n1_adj_220), .I0(state[7]), .I1(n5984));
    AND2 select_163_Select_66_i2 (.O(n2_adj_49), .I0(state[6]), .I1(dataInBuf[58]));
    OR3 i1_adj_5 (.O(n5683), .I0(n2_adj_304), .I1(n1_adj_303), .I2(state[0]));
    AND2 select_163_Select_65_i2 (.O(n2_adj_47), .I0(state[6]), .I1(dataInBuf[57]));
    OR2 select_163_Select_64_i9 (.O(n9_adj_45), .I0(n2_adj_44), .I1(n1_adj_43));
    AND2 select_163_Select_142_i1 (.O(n1_adj_217), .I0(state[7]), .I1(n5981));
    AND2 select_163_Select_64_i2 (.O(n2_adj_44), .I0(state[6]), .I1(dataInBuf[56]));
    AND2 select_163_Select_141_i1 (.O(n1_adj_215), .I0(state[7]), .I1(n5978));
    AND2 select_163_Select_140_i1 (.O(n1_adj_212), .I0(state[7]), .I1(n5975));
    AND2 select_163_Select_139_i1 (.O(n1_adj_209), .I0(state[7]), .I1(n5972));
    AND2 select_163_Select_138_i1 (.O(n1_adj_206), .I0(state[7]), .I1(n5969));
    AND2 select_163_Select_62_i2 (.O(n2_adj_42), .I0(state[6]), .I1(dataInBuf[54]));
    OR2 select_163_Select_61_i9 (.O(n9_adj_40), .I0(n2_adj_39), .I1(n1_adj_38));
    AND2 select_163_Select_61_i2 (.O(n2_adj_39), .I0(state[6]), .I1(dataInBuf[53]));
    AND2 select_163_Select_137_i1 (.O(n1_adj_203), .I0(state[7]), .I1(n5966));
    XOR2 i2301 (.O(n94), .I0(n5120), .I1(cnt[11]));
    OR2 select_163_Select_58_i9 (.O(n9_adj_37), .I0(n2_adj_36), .I1(n1_adj_35));
    AND2 select_163_Select_58_i2 (.O(n2_adj_36), .I0(state[6]), .I1(dataInBuf[50]));
    AND2 select_163_Select_136_i1 (.O(n1_adj_200), .I0(state[7]), .I1(n5963));
    OR2 i3202 (.O(n6023), .I0(n6022), .I1(n6021));
    OR3 i2_adj_6 (.O(n5255), .I0(n1_adj_7), .I1(state[0]), .I2(n2_adj_8));
    AND2 select_163_Select_134_i1 (.O(n1_adj_197), .I0(state[7]), .I1(n5960));
    AND2 select_163_Select_57_i2 (.O(n2_adj_34), .I0(state[6]), .I1(dataInBuf[49]));
    OR2 i3139 (.O(n5960), .I0(n5959), .I1(n5958));
    AND2 select_163_Select_56_i2 (.O(n2_adj_32), .I0(state[6]), .I1(dataInBuf[48]));
    AND2 i2290 (.O(n5113), .I0(n5106), .I1(cnt[9]));
    AND2 select_163_Select_133_i1 (.O(n1_adj_195), .I0(state[7]), .I1(n5957));
    AND2 select_163_Select_132_i1 (.O(n1_adj_192), .I0(state[7]), .I1(n5954));
    AND2 select_163_Select_54_i2 (.O(n2_adj_30), .I0(state[6]), .I1(dataInBuf[46]));
    OR2 select_163_Select_53_i9 (.O(n9_adj_28), .I0(n2_adj_27), .I1(n1_adj_26));
    AND2 select_163_Select_131_i1 (.O(n1_adj_189), .I0(state[7]), .I1(n5951));
    AND2 select_163_Select_130_i1 (.O(n1_adj_186), .I0(state[7]), .I1(n5948));
    AND2 select_163_Select_53_i2 (.O(n2_adj_27), .I0(state[6]), .I1(dataInBuf[45]));
    AND2 select_163_Select_129_i1 (.O(n1_adj_183), .I0(state[7]), .I1(n5945));
    AND2 select_163_Select_128_i1 (.O(n1_adj_180), .I0(state[7]), .I1(n5942));
    AND2 select_163_Select_126_i1 (.O(n1_adj_177), .I0(state[7]), .I1(n5939));
    AND2 i3141 (.O(n5962), .I0(lcdRs_N_619), .I1(dataInBuf[136]));
    AND2 select_163_Select_125_i1 (.O(n1_adj_175), .I0(state[7]), .I1(n5936));
    XOR2 i2308 (.O(n93), .I0(n5127), .I1(cnt[12]));
    XOR2 i2238 (.O(n103), .I0(n5057), .I1(cnt[2]));
    OR2 select_162_Select_0_i9 (.O(lcdRs_N_615), .I0(state[6]), .I1(n1_adj_25));
    AND2 select_163_Select_124_i1 (.O(n1_adj_172), .I0(state[7]), .I1(n5933));
    AND2 select_163_Select_123_i1 (.O(n1_adj_169), .I0(state[7]), .I1(n5930));
    AND2 select_163_Select_122_i1 (.O(n1_adj_166), .I0(state[7]), .I1(n5927));
    AND2 i3228 (.O(n6049), .I0(lcdRs_N_619), .I1(dataInBuf[169]));
    OR2 i2907 (.O(n5729), .I0(state[4]), .I1(n20));
    OR2 i2920 (.O(n5741), .I0(n5740), .I1(n5739));
    OR2 i3229 (.O(n6050), .I0(n6049), .I1(n6048));
    AND2 i3231 (.O(n6052), .I0(lcdRs_N_619), .I1(dataInBuf[170]));
    OR2 i3232 (.O(n6053), .I0(n6052), .I1(n6051));
    OR4 i3 (.O(n5258), .I0(n3012), .I1(state[4]), .I2(n20), .I3(state[1]));
    AND2 i3234 (.O(n6055), .I0(lcdRs_N_619), .I1(dataInBuf[171]));
    OR2 i3235 (.O(n6056), .I0(n6055), .I1(n6054));
    AND2 i3237 (.O(n6058), .I0(lcdRs_N_619), .I1(dataInBuf[172]));
    OR2 i3238 (.O(n6059), .I0(n6058), .I1(n6057));
    AND2 i2917 (.O(n3804), .I0(n5737), .I1(n1_adj_482));
    AND2 i3240 (.O(n6061), .I0(lcdRs_N_619), .I1(dataInBuf[173]));
    OR2 i3241 (.O(n6062), .I0(n6061), .I1(n6060));
    OR2 i2926 (.O(n5747), .I0(n5746), .I1(n5745));
    AND2 i3243 (.O(n6064), .I0(lcdRs_N_619), .I1(dataInBuf[174]));
    OR2 i3244 (.O(n6065), .I0(n6064), .I1(n6063));
    AND2 i2928 (.O(n5749), .I0(lcdRs_N_619), .I1(dataInBuf[37]));
    AND2 i3246 (.O(n6067), .I0(lcdRs_N_619), .I1(dataInBuf[176]));
    OR2 i3247 (.O(n6068), .I0(n6067), .I1(n6066));
    OR2 i2929 (.O(n5750), .I0(n5749), .I1(n5748));
    AND2 i3249 (.O(n6070), .I0(lcdRs_N_619), .I1(dataInBuf[177]));
    OR2 i3250 (.O(n6071), .I0(n6070), .I1(n6069));
    AND2 i2931 (.O(n5752), .I0(lcdRs_N_619), .I1(dataInBuf[41]));
    AND2 i3252 (.O(n6073), .I0(lcdRs_N_619), .I1(dataInBuf[178]));
    OR2 i3253 (.O(n6074), .I0(n6073), .I1(n6072));
    OR2 i2932 (.O(n5753), .I0(n5752), .I1(n5751));
    AND2 i3255 (.O(n6076), .I0(lcdRs_N_619), .I1(dataInBuf[179]));
    OR2 i3256 (.O(n6077), .I0(n6076), .I1(n6075));
    AND2 i2934 (.O(n5755), .I0(lcdRs_N_619), .I1(dataInBuf[42]));
    AND2 i3258 (.O(n6079), .I0(lcdRs_N_619), .I1(dataInBuf[180]));
    OR2 i3259 (.O(n6080), .I0(n6079), .I1(n6078));
    OR2 i2935 (.O(n5756), .I0(n5755), .I1(n5754));
    AND2 i3261 (.O(n6082), .I0(lcdRs_N_619), .I1(dataInBuf[181]));
    OR2 i3262 (.O(n6083), .I0(n6082), .I1(n6081));
    AND2 i2937 (.O(n5758), .I0(lcdRs_N_619), .I1(dataInBuf[45]));
    OR2 select_163_Select_45_i9 (.O(n9_adj_24), .I0(n2_adj_23), .I1(n1_adj_22));
    AND2 i3264 (.O(n6085), .I0(lcdRs_N_619), .I1(dataInBuf[182]));
    OR2 i3265 (.O(n6086), .I0(n6085), .I1(n6084));
    OR2 i2938 (.O(n5759), .I0(n5758), .I1(n5757));
    AND2 i2918 (.O(n5739), .I0(lcdRs_N_618), .I1(dataInBuf[5]));
    AND2 i3267 (.O(n6088), .I0(lcdRs_N_619), .I1(dataInBuf[184]));
    OR2 i3268 (.O(n6089), .I0(n6088), .I1(n6087));
    AND2 select_163_Select_121_i1 (.O(n1_adj_163), .I0(state[7]), .I1(n5924));
    AND2 i2940 (.O(n5761), .I0(lcdRs_N_619), .I1(dataInBuf[46]));
    OR2 i2941 (.O(n5762), .I0(n5761), .I1(n5760));
    AND2 i3270 (.O(n6091), .I0(lcdRs_N_619), .I1(dataInBuf[185]));
    OR2 i1_adj_7 (.O(n7), .I0(n5734), .I1(n3800));
    OR2 i3271 (.O(n6092), .I0(n6091), .I1(n6090));
    AND2 i1_adj_8 (.O(n5650), .I0(n7), .I1(state[7]));
    OR3 i1_adj_9 (.O(n5693), .I0(n2_adj_176), .I1(n1_adj_175), .I2(state[0]));
    OR2 select_163_Select_254_i9 (.O(n9_adj_481), .I0(n2_adj_480), .I1(n1_adj_479));
    OR3 i1_adj_10 (.O(n5661), .I0(n1_adj_11), .I1(n2_adj_12), .I2(state[0]));
    AND2 i3273 (.O(n6094), .I0(lcdRs_N_619), .I1(dataInBuf[186]));
    OR3 i1_adj_11 (.O(n5663), .I0(n1_adj_20), .I1(n2_adj_21), .I2(state[0]));
    AND2 i2943 (.O(n5764), .I0(lcdRs_N_619), .I1(dataInBuf[49]));
    AND2 select_163_Select_254_i2 (.O(n2_adj_480), .I0(state[6]), .I1(dataInBuf[246]));
    OR2 i3274 (.O(n6095), .I0(n6094), .I1(n6093));
    AND2 i3276 (.O(n6097), .I0(lcdRs_N_619), .I1(dataInBuf[187]));
    OR3 i1_adj_12 (.O(n5659), .I0(n2_adj_456), .I1(n1_adj_455), .I2(state[0]));
    OR2 i2944 (.O(n5765), .I0(n5764), .I1(n5763));
    OR3 i1_adj_13 (.O(n5695), .I0(n2_adj_96), .I1(n1_adj_95), .I2(state[0]));
    AND2 select_163_Select_253_i2 (.O(n2_adj_478), .I0(state[6]), .I1(dataInBuf[245]));
    OR3 i1_adj_14 (.O(n5697), .I0(n2_adj_70), .I1(n1_adj_69), .I2(state[0]));
    OR2 i3277 (.O(n6098), .I0(n6097), .I1(n6096));
    AND2 i2946 (.O(n5767), .I0(lcdRs_N_619), .I1(dataInBuf[50]));
    OR2 select_163_Select_252_i9 (.O(n9_adj_476), .I0(n2_adj_475), .I1(n1_adj_474));
    OR2 i2947 (.O(n5768), .I0(n5767), .I1(n5766));
    AND2 select_163_Select_252_i2 (.O(n2_adj_475), .I0(state[6]), .I1(dataInBuf[244]));
    OR2 select_163_Select_251_i9 (.O(n9_adj_473), .I0(n2_adj_472), .I1(n1_adj_471));
    AND2 select_163_Select_251_i2 (.O(n2_adj_472), .I0(state[6]), .I1(dataInBuf[243]));
    OR2 select_163_Select_250_i9 (.O(n9_adj_470), .I0(n2_adj_469), .I1(n1_adj_468));
    AND2 select_163_Select_250_i2 (.O(n2_adj_469), .I0(state[6]), .I1(dataInBuf[242]));
    OR2 select_163_Select_249_i9 (.O(n9_adj_467), .I0(n2_adj_466), .I1(n1_adj_465));
    AND2 select_163_Select_249_i2 (.O(n2_adj_466), .I0(state[6]), .I1(dataInBuf[241]));
    OR2 select_163_Select_248_i9 (.O(n9_adj_464), .I0(n2_adj_463), .I1(n1_adj_462));
    AND2 select_163_Select_248_i2 (.O(n2_adj_463), .I0(state[6]), .I1(dataInBuf[240]));
    XOR2 i2231 (.O(n104), .I0(cnt[0]), .I1(cnt[1]));
    OR2 select_163_Select_246_i9 (.O(n9_adj_459), .I0(n2_adj_458), .I1(n1_adj_457));
    AND2 select_163_Select_246_i2 (.O(n2_adj_458), .I0(state[6]), .I1(dataInBuf[238]));
    AND2 select_163_Select_245_i2 (.O(n2_adj_456), .I0(state[6]), .I1(dataInBuf[237]));
    OR2 select_163_Select_244_i9 (.O(n9_adj_454), .I0(n2_adj_453), .I1(n1_adj_452));
    AND2 select_163_Select_244_i2 (.O(n2_adj_453), .I0(state[6]), .I1(dataInBuf[236]));
    OR2 select_163_Select_243_i9 (.O(n9_adj_451), .I0(n2_adj_450), .I1(n1_adj_449));
    AND2 select_163_Select_243_i2 (.O(n2_adj_450), .I0(state[6]), .I1(dataInBuf[235]));
    OR2 select_163_Select_242_i9 (.O(n9_adj_448), .I0(n2_adj_447), .I1(n1_adj_446));
    AND2 select_163_Select_242_i2 (.O(n2_adj_447), .I0(state[6]), .I1(dataInBuf[234]));
    OR2 select_163_Select_241_i9 (.O(n9_adj_445), .I0(n2_adj_444), .I1(n1_adj_443));
    AND2 select_163_Select_241_i2 (.O(n2_adj_444), .I0(state[6]), .I1(dataInBuf[233]));
    OR2 select_163_Select_240_i9 (.O(n9_adj_442), .I0(n2_adj_441), .I1(n1_adj_440));
    AND2 select_163_Select_240_i2 (.O(n2_adj_441), .I0(state[6]), .I1(dataInBuf[232]));
    AND2 i2255 (.O(n5078), .I0(n5071), .I1(cnt[4]));
    OR2 select_163_Select_238_i9 (.O(n9_adj_439), .I0(n2_adj_438), .I1(n1_adj_437));
    AND2 select_163_Select_238_i2 (.O(n2_adj_438), .I0(state[6]), .I1(dataInBuf[230]));
    OR2 i2_adj_15 (.O(n3649), .I0(n1_adj_482), .I1(state[0]));
    AND2 select_163_Select_237_i2 (.O(n2_adj_436), .I0(state[6]), .I1(dataInBuf[229]));
    OR2 select_163_Select_236_i9 (.O(n9_adj_434), .I0(n2_adj_433), .I1(n1_adj_432));
    AND2 i2949 (.O(n5770), .I0(lcdRs_N_619), .I1(dataInBuf[53]));
    OR2 select_105_i5 (.O(n20), .I0(state[3]), .I1(state[2]));
    AND2 select_163_Select_236_i2 (.O(n2_adj_433), .I0(state[6]), .I1(dataInBuf[228]));
    AND2 i3279 (.O(n6100), .I0(lcdRs_N_619), .I1(dataInBuf[188]));
    OR2 i2950 (.O(n5771), .I0(n5770), .I1(n5769));
    OR2 select_105_i9 (.O(n40), .I0(n2185), .I1(n3012));
    OR2 select_163_Select_235_i9 (.O(n9_adj_431), .I0(n2_adj_430), .I1(n1_adj_429));
    AND2 select_163_Select_45_i2 (.O(n2_adj_23), .I0(state[6]), .I1(dataInBuf[37]));
    OR2 i3280 (.O(n6101), .I0(n6100), .I1(n6099));
    OR2 select_105_i13 (.O(n60), .I0(n40), .I1(state[4]));
    AND2 i3282 (.O(n6103), .I0(lcdRs_N_619), .I1(dataInBuf[189]));
    AND2 select_163_Select_120_i1 (.O(n1_adj_160), .I0(state[7]), .I1(n5921));
    AND2 i2952 (.O(n5773), .I0(lcdRs_N_619), .I1(dataInBuf[54]));
    AND2 select_163_Select_235_i2 (.O(n2_adj_430), .I0(state[6]), .I1(dataInBuf[227]));
    OR2 i3283 (.O(n6104), .I0(n6103), .I1(n6102));
    AND2 i3285 (.O(n6106), .I0(lcdRs_N_619), .I1(dataInBuf[190]));
    OR2 select_163_Select_234_i9 (.O(n9_adj_428), .I0(n2_adj_427), .I1(n1_adj_426));
    OR2 i2953 (.O(n5774), .I0(n5773), .I1(n5772));
    OR2 i3286 (.O(n6107), .I0(n6106), .I1(n6105));
    AND2 i3288 (.O(n6109), .I0(lcdRs_N_619), .I1(dataInBuf[192]));
    AND2 i2955 (.O(n5776), .I0(lcdRs_N_619), .I1(dataInBuf[56]));
    AND2 select_163_Select_234_i2 (.O(n2_adj_427), .I0(state[6]), .I1(dataInBuf[226]));
    OR2 i3289 (.O(n6110), .I0(n6109), .I1(n6108));
    OR2 select_163_Select_233_i9 (.O(n9_adj_425), .I0(n2_adj_424), .I1(n1_adj_423));
    AND2 select_163_Select_233_i2 (.O(n2_adj_424), .I0(state[6]), .I1(dataInBuf[225]));
    OR2 select_163_Select_232_i9 (.O(n9_adj_422), .I0(n2_adj_421), .I1(n1_adj_420));
    AND2 select_163_Select_232_i2 (.O(n2_adj_421), .I0(state[6]), .I1(dataInBuf[224]));
    AND2 i2339 (.O(n5162), .I0(n5155), .I1(cnt[16]));
    OR2 select_163_Select_230_i9 (.O(n9_adj_419), .I0(n2_adj_418), .I1(n1_adj_417));
    AND2 select_163_Select_230_i2 (.O(n2_adj_418), .I0(state[6]), .I1(dataInBuf[222]));
    AND2 i3291 (.O(n6112), .I0(lcdRs_N_619), .I1(dataInBuf[193]));
    OR3 i1_adj_16 (.O(n5699), .I0(n2_adj_47), .I1(n1_adj_46), .I2(state[0]));
    AND2 select_163_Select_229_i2 (.O(n2_adj_416), .I0(state[6]), .I1(dataInBuf[221]));
    OR2 select_163_Select_228_i9 (.O(n9_adj_414), .I0(n2_adj_413), .I1(n1_adj_412));
    AND2 select_163_Select_228_i2 (.O(n2_adj_413), .I0(state[6]), .I1(dataInBuf[220]));
    OR2 select_163_Select_227_i9 (.O(n9_adj_411), .I0(n2_adj_410), .I1(n1_adj_409));
    AND2 select_163_Select_227_i2 (.O(n2_adj_410), .I0(state[6]), .I1(dataInBuf[219]));
    OR2 select_163_Select_226_i9 (.O(n9_adj_408), .I0(n2_adj_407), .I1(n1_adj_406));
    AND2 select_163_Select_226_i2 (.O(n2_adj_407), .I0(state[6]), .I1(dataInBuf[218]));
    OR2 select_163_Select_225_i9 (.O(n9_adj_405), .I0(n2_adj_404), .I1(n1_adj_403));
    AND2 select_163_Select_225_i2 (.O(n2_adj_404), .I0(state[6]), .I1(dataInBuf[217]));
    OR2 select_163_Select_224_i9 (.O(n9_adj_402), .I0(n2_adj_401), .I1(n1_adj_400));
    AND2 select_163_Select_224_i2 (.O(n2_adj_401), .I0(state[6]), .I1(dataInBuf[216]));
    OR2 select_163_Select_222_i9 (.O(n9_adj_399), .I0(n2_adj_398), .I1(n1_adj_397));
    AND2 select_163_Select_222_i2 (.O(n2_adj_398), .I0(state[6]), .I1(dataInBuf[214]));
    AND2 select_163_Select_221_i2 (.O(n2_adj_396), .I0(state[6]), .I1(dataInBuf[213]));
    AND2 select_163_Select_220_i2 (.O(n2_adj_394), .I0(state[6]), .I1(dataInBuf[212]));
    OR2 select_163_Select_219_i9 (.O(n9_adj_392), .I0(n2_adj_391), .I1(n1_adj_390));
    AND2 select_163_Select_219_i2 (.O(n2_adj_391), .I0(state[6]), .I1(dataInBuf[211]));
    AND2 i3461 (.O(n6282), .I0(n4374), .I1(n3100));
    AND2 i1550 (.O(n3638), .I0(n4374), .I1(n3637));
    OR3 i1_adj_17 (.O(n5691), .I0(n2_adj_236), .I1(n1_adj_235), .I2(state[0]));
    AND2 select_163_Select_118_i1 (.O(n1_adj_157), .I0(state[7]), .I1(n5918));
    AND2 select_163_Select_117_i1 (.O(n1_adj_155), .I0(state[7]), .I1(n5915));
    OR2 i3142 (.O(n5963), .I0(n5962), .I1(n5961));
    AND2 select_163_Select_46_i2 (.O(n2_adj_21), .I0(state[6]), .I1(dataInBuf[38]));
    AND2 i2297 (.O(n5120), .I0(n5113), .I1(cnt[10]));
    XOR2 i2315 (.O(n92), .I0(n5134), .I1(cnt[13]));
    AND2 select_163_Select_116_i1 (.O(n1_adj_152), .I0(state[7]), .I1(n5912));
    AND2 select_163_Select_115_i1 (.O(n1_adj_149), .I0(state[7]), .I1(n5909));
    AND2 select_163_Select_114_i1 (.O(n1_adj_146), .I0(state[7]), .I1(n5906));
    AND2 i3144 (.O(n5965), .I0(lcdRs_N_619), .I1(dataInBuf[137]));
    OR2 i3145 (.O(n5966), .I0(n5965), .I1(n5964));
    AND2 i3147 (.O(n5968), .I0(lcdRs_N_619), .I1(dataInBuf[138]));
    AND2 select_163_Select_113_i1 (.O(n1_adj_143), .I0(state[7]), .I1(n5903));
    OR2 select_163_Select_5_i13 (.O(n3000), .I0(state[0]), .I1(n5724));
    AND2 select_163_Select_112_i1 (.O(n1_adj_140), .I0(state[7]), .I1(n5900));
    AND2 select_163_Select_110_i1 (.O(n1_adj_137), .I0(state[7]), .I1(n5897));
    AND2 select_163_Select_109_i1 (.O(n1_adj_135), .I0(state[7]), .I1(n5894));
    OR2 i3148 (.O(n5969), .I0(n5968), .I1(n5967));
    OR3 i2_adj_18 (.O(n5259), .I0(n1_adj_1), .I1(state[0]), .I2(n2));
    AND2 select_163_Select_108_i1 (.O(n1_adj_132), .I0(state[7]), .I1(n5891));
    AND2 select_163_Select_107_i1 (.O(n1_adj_129), .I0(state[7]), .I1(n5888));
    AND2 select_163_Select_13_i2 (.O(n2_adj_19), .I0(state[6]), .I1(dataInBuf[5]));
    AND2 i3150 (.O(n5971), .I0(lcdRs_N_619), .I1(dataInBuf[139]));
    OR2 i3151 (.O(n5972), .I0(n5971), .I1(n5970));
    AND2 select_163_Select_106_i1 (.O(n1_adj_126), .I0(state[7]), .I1(n5885));
    AND2 select_163_Select_105_i1 (.O(n1_adj_123), .I0(state[7]), .I1(n5882));
    AND2 select_163_Select_104_i1 (.O(n1_adj_120), .I0(state[7]), .I1(n5879));
    AND2 i3153 (.O(n5974), .I0(lcdRs_N_619), .I1(dataInBuf[140]));
    AND2 select_163_Select_102_i1 (.O(n1_adj_117), .I0(state[7]), .I1(n5876));
    OR3 i1_adj_19 (.O(n5685), .I0(n2_adj_289), .I1(n1_adj_288), .I2(state[0]));
    AND2 select_163_Select_101_i1 (.O(n1_adj_115), .I0(state[7]), .I1(n5873));
    AND2 i2248 (.O(n5071), .I0(n5064), .I1(cnt[3]));
    OR2 i3154 (.O(n5975), .I0(n5974), .I1(n5973));
    AND2 i3156 (.O(n5977), .I0(lcdRs_N_619), .I1(dataInBuf[141]));
    AND2 select_163_Select_100_i1 (.O(n1_adj_112), .I0(state[7]), .I1(n5870));
    OR2 select_163_Select_37_i9 (.O(n9_adj_17), .I0(n2_adj_16), .I1(n1_adj_15));
    AND2 select_163_Select_99_i1 (.O(n1_adj_109), .I0(state[7]), .I1(n5867));
    AND2 select_163_Select_98_i1 (.O(n1_adj_106), .I0(state[7]), .I1(n5864));
    AND2 select_163_Select_37_i2 (.O(n2_adj_16), .I0(state[6]), .I1(dataInBuf[29]));
    OR2 i3157 (.O(n5978), .I0(n5977), .I1(n5976));
    AND2 i3159 (.O(n5980), .I0(lcdRs_N_619), .I1(dataInBuf[142]));
    AND2 select_163_Select_97_i1 (.O(n1_adj_103), .I0(state[7]), .I1(n5861));
    AND2 select_163_Select_96_i1 (.O(n1_adj_100), .I0(state[7]), .I1(n5858));
    AND2 select_163_Select_94_i1 (.O(n1_adj_97), .I0(state[7]), .I1(n5855));
    AND2 select_163_Select_93_i1 (.O(n1_adj_95), .I0(state[7]), .I1(n5852));
    AND2 select_163_Select_92_i1 (.O(n1_adj_93), .I0(state[7]), .I1(n5849));
    OR2 select_163_Select_49_i9 (.O(n9_adj_14), .I0(n2_adj_4), .I1(n1_adj_5));
    AND2 select_163_Select_49_i2 (.O(n2_adj_4), .I0(state[6]), .I1(dataInBuf[41]));
    OR2 i1_adj_20 (.O(n4_adj_460), .I0(state[0]), .I1(n5727));
    AND2 select_163_Select_91_i1 (.O(n1_adj_91), .I0(state[7]), .I1(n5846));
    AND2 select_163_Select_90_i1 (.O(n1_adj_88), .I0(state[7]), .I1(n5843));
    AND2 select_163_Select_89_i1 (.O(n1_adj_85), .I0(state[7]), .I1(n5840));
    AND2 select_163_Select_88_i1 (.O(n1_adj_82), .I0(state[7]), .I1(n5837));
    AND2 i3204 (.O(n6025), .I0(lcdRs_N_619), .I1(dataInBuf[160]));
    AND2 select_163_Select_50_i2 (.O(n2_adj_8), .I0(state[6]), .I1(dataInBuf[42]));
    OR2 i3160 (.O(n5981), .I0(n5980), .I1(n5979));
    OR2 select_163_Select_41_i9 (.O(n9), .I0(n2_adj_13), .I1(n1_adj_9));
    AND2 select_163_Select_41_i2 (.O(n2_adj_13), .I0(state[6]), .I1(dataInBuf[33]));
    AND2 select_163_Select_86_i1 (.O(n1_adj_79), .I0(state[7]), .I1(n5834));
    XOR2 i2322 (.O(n91), .I0(n5141), .I1(cnt[14]));
    AND2 select_163_Select_85_i1 (.O(n1_adj_77), .I0(state[7]), .I1(n5831));
    AND2 i2304 (.O(n5127), .I0(n5120), .I1(cnt[11]));
    AND2 select_163_Select_42_i2 (.O(n2_adj_3), .I0(state[6]), .I1(dataInBuf[34]));
    AND2 select_163_Select_82_i1 (.O(n1_adj_74), .I0(state[7]), .I1(n5828));
    AND2 select_163_Select_81_i1 (.O(n1_adj_71), .I0(state[7]), .I1(n5825));
    OR2 i1_adj_21 (.O(n4_adj_461), .I0(state[0]), .I1(n5725));
    AND2 select_163_Select_29_i2 (.O(n2), .I0(state[6]), .I1(dataInBuf[21]));
    AND2 select_163_Select_80_i1 (.O(n1_adj_69), .I0(state[7]), .I1(n5822));
    AND2 select_163_Select_78_i1 (.O(n1_adj_67), .I0(state[7]), .I1(n5819));
    AND2 select_163_Select_77_i1 (.O(n1_adj_64), .I0(state[7]), .I1(n5816));
    XOR2 i2245 (.O(n102), .I0(n5064), .I1(cnt[3]));
    AND2 i3162 (.O(n5983), .I0(lcdRs_N_619), .I1(dataInBuf[144]));
    AND2 select_163_Select_74_i1 (.O(n1_adj_61), .I0(state[7]), .I1(n5813));
    AND2 select_163_Select_21_i2 (.O(n2_adj_12), .I0(state[6]), .I1(dataInBuf[13]));
    AND2 select_163_Select_73_i1 (.O(n1_adj_58), .I0(state[7]), .I1(n5810));
    OR3 i2_adj_22 (.O(n5196), .I0(n1_adj_215), .I1(n2_adj_216), .I2(state[0]));
    AND2 select_163_Select_72_i1 (.O(n1_adj_56), .I0(state[7]), .I1(n5807));
    AND2 select_163_Select_70_i1 (.O(n1_adj_54), .I0(state[7]), .I1(n5804));
    OR2 i3163 (.O(n5984), .I0(n5983), .I1(n5982));
    AND2 select_163_Select_69_i1 (.O(n1_adj_51), .I0(state[7]), .I1(n5801));
    AND2 i3165 (.O(n5986), .I0(lcdRs_N_619), .I1(dataInBuf[145]));
    OR2 i3166 (.O(n5987), .I0(n5986), .I1(n5985));
    AND2 i3168 (.O(n5989), .I0(lcdRs_N_619), .I1(dataInBuf[146]));
    OR2 i3205 (.O(n6026), .I0(n6025), .I1(n6024));
    OR2 i3169 (.O(n5990), .I0(n5989), .I1(n5988));
    AND2 i3207 (.O(n6028), .I0(lcdRs_N_619), .I1(dataInBuf[161]));
    AND2 select_163_Select_66_i1 (.O(n1_adj_48), .I0(state[7]), .I1(n5798));
    AND2 i3171 (.O(n5992), .I0(lcdRs_N_619), .I1(dataInBuf[147]));
    AND2 select_163_Select_65_i1 (.O(n1_adj_46), .I0(state[7]), .I1(n5795));
    XOR2 i2329 (.O(n90), .I0(n5148), .I1(cnt[15]));
    OR2 i3172 (.O(n5993), .I0(n5992), .I1(n5991));
    OR3 i1_adj_23 (.O(n5687), .I0(n2_adj_272), .I1(n1_adj_271), .I2(state[0]));
    AND2 select_163_Select_64_i1 (.O(n1_adj_43), .I0(state[7]), .I1(n5792));
    AND6 i19 (.O(n5194), .I0(n36), .I1(cnt[13]), .I2(n26), .I3(n34), 
         .I4(n35), .I5(cnt[8]));
    AND2 select_163_Select_62_i1 (.O(n1_adj_41), .I0(state[7]), .I1(n5789));
    OR3 i2_adj_24 (.O(n5218), .I0(n1_adj_305), .I1(n2_adj_306), .I2(state[0]));
    AND2 i3174 (.O(n5995), .I0(lcdRs_N_619), .I1(dataInBuf[148]));
    OR2 i3175 (.O(n5996), .I0(n5995), .I1(n5994));
    XOR2 i202 (.O(dispCount_5__N_347[2]), .I0(n3033), .I1(dispCount[2]));
    AND2 i218 (.O(n3054), .I0(n3047), .I1(dispCount[4]));
    AND2 select_163_Select_61_i1 (.O(n1_adj_38), .I0(state[7]), .I1(n5786));
    OR2 i3208 (.O(n6029), .I0(n6028), .I1(n6027));
    AND2 i204 (.O(n3040), .I0(n3033), .I1(dispCount[2]));
    AND2 select_163_Select_58_i1 (.O(n1_adj_35), .I0(state[7]), .I1(n5783));
    AND2 i197 (.O(n3033), .I0(dispCount[0]), .I1(dispCount[1]));
    AND2 select_163_Select_57_i1 (.O(n1_adj_33), .I0(state[7]), .I1(n5780));
    AND2 i211 (.O(n3047), .I0(n3040), .I1(dispCount[3]));
    XOR2 i195 (.O(dispCount_5__N_347[1]), .I0(dispCount[0]), .I1(dispCount[1]));
    AND2 select_163_Select_56_i1 (.O(n1_adj_31), .I0(state[7]), .I1(n5777));
    AND2 select_163_Select_54_i1 (.O(n1_adj_29), .I0(state[7]), .I1(n5774));
    OR2 i1_adj_25 (.O(n14), .I0(n3731), .I1(n1));
    AND2 select_163_Select_53_i1 (.O(n1_adj_26), .I0(state[7]), .I1(n5771));
    AND2 i1_adj_26 (.O(n2212), .I0(lcdRs_N_620), .I1(state[7]));
    XOR2 i216 (.O(dispCount_5__N_347[4]), .I0(n3047), .I1(dispCount[4]));
    AND2 i3210 (.O(n6031), .I0(lcdRs_N_619), .I1(dataInBuf[162]));
    XOR2 i223 (.O(dispCount_5__N_347[5]), .I0(n3054), .I1(dispCount[5]));
    AND2 i3177 (.O(n5998), .I0(lcdRs_N_619), .I1(dataInBuf[149]));
    AND2 select_162_Select_0_i1 (.O(n1_adj_25), .I0(state[7]), .I1(lcdRs_N_617));
    OR2 i3178 (.O(n5999), .I0(n5998), .I1(n5997));
    OR2 i3211 (.O(n6032), .I0(n6031), .I1(n6030));
    AND2 i2925 (.O(n5746), .I0(lcdRs_N_619), .I1(dataInBuf[29]));
    XOR2 i32 (.O(n16), .I0(dispCount[5]), .I1(dispCount[4]));
    AND2 select_163_Select_45_i1 (.O(n1_adj_22), .I0(state[7]), .I1(n5759));
    AND3 i3455 (.O(n6276), .I0(n4376), .I1(n4374), .I2(n3117));
    AND2 i3452 (.O(n6273), .I0(lcdRs_N_618), .I1(dataInBuf[246]));
    AND2 i3449 (.O(n6270), .I0(lcdRs_N_618), .I1(dataInBuf[245]));
    AND2 select_163_Select_46_i1 (.O(n1_adj_20), .I0(state[7]), .I1(n5762));
    OR3 i2_adj_27 (.O(n5210), .I0(n1_adj_415), .I1(n2_adj_416), .I2(state[0]));
    AND2 i3213 (.O(n6034), .I0(lcdRs_N_619), .I1(dataInBuf[163]));
    OR2 reduce_or_136_i1 (.O(n2185), .I0(n3006), .I1(state[6]));
    AND2 i3446 (.O(n6267), .I0(lcdRs_N_618), .I1(dataInBuf[244]));
    AND2 i3443 (.O(n6264), .I0(lcdRs_N_618), .I1(dataInBuf[243]));
    AND2 i3440 (.O(n6261), .I0(lcdRs_N_618), .I1(dataInBuf[242]));
    AND2 i3437 (.O(n6258), .I0(lcdRs_N_618), .I1(dataInBuf[241]));
    OR2 i3214 (.O(n6035), .I0(n6034), .I1(n6033));
    AND2 i3216 (.O(n6037), .I0(lcdRs_N_619), .I1(dataInBuf[164]));
    OR2 i3217 (.O(n6038), .I0(n6037), .I1(n6036));
    AND2 i3219 (.O(n6040), .I0(lcdRs_N_619), .I1(dataInBuf[165]));
    XOR2 i2336 (.O(n89), .I0(n5155), .I1(cnt[16]));
    AND2 i3434 (.O(n6255), .I0(lcdRs_N_618), .I1(dataInBuf[240]));
    AND2 i3431 (.O(n6252), .I0(lcdRs_N_618), .I1(dataInBuf[238]));
    AND2 i2241 (.O(n5064), .I0(n5057), .I1(cnt[2]));
    AND2 i3428 (.O(n6249), .I0(lcdRs_N_618), .I1(dataInBuf[237]));
    OR2 i1_adj_28 (.O(n3733), .I0(n5721), .I1(state[0]));
    OR2 i3220 (.O(n6041), .I0(n6040), .I1(n6039));
    AND2 i3222 (.O(n6043), .I0(lcdRs_N_619), .I1(dataInBuf[166]));
    AND2 i3425 (.O(n6246), .I0(lcdRs_N_618), .I1(dataInBuf[236]));
    AND2 select_163_Select_13_i1 (.O(n1_adj_18), .I0(state[7]), .I1(n5741));
    AND2 i3422 (.O(n6243), .I0(lcdRs_N_618), .I1(dataInBuf[235]));
    AND2 i3419 (.O(n6240), .I0(lcdRs_N_618), .I1(dataInBuf[234]));
    OR2 i3223 (.O(n6044), .I0(n6043), .I1(n6042));
    AND2 i3416 (.O(n6237), .I0(lcdRs_N_618), .I1(dataInBuf[233]));
    AND2 select_163_Select_37_i1 (.O(n1_adj_15), .I0(state[7]), .I1(n5750));
    AND2 i3225 (.O(n6046), .I0(lcdRs_N_619), .I1(dataInBuf[168]));
    AND2 i3413 (.O(n6234), .I0(lcdRs_N_618), .I1(dataInBuf[232]));
    AND2 select_163_Select_49_i1 (.O(n1_adj_5), .I0(state[7]), .I1(n5765));
    AND2 i3410 (.O(n6231), .I0(lcdRs_N_618), .I1(dataInBuf[230]));
    AND2 select_163_Select_50_i1 (.O(n1_adj_7), .I0(state[7]), .I1(n5768));
    AND2 i3407 (.O(n6228), .I0(lcdRs_N_618), .I1(dataInBuf[229]));
    AND2 i3404 (.O(n6225), .I0(lcdRs_N_618), .I1(dataInBuf[228]));
    AND2 i3401 (.O(n6222), .I0(lcdRs_N_618), .I1(dataInBuf[227]));
    AND2 select_163_Select_41_i1 (.O(n1_adj_9), .I0(state[7]), .I1(n5753));
    AND2 i3398 (.O(n6219), .I0(lcdRs_N_618), .I1(dataInBuf[226]));
    AND2 select_163_Select_42_i1 (.O(n1_adj_2), .I0(state[7]), .I1(n5756));
    AND2 i3395 (.O(n6216), .I0(lcdRs_N_618), .I1(dataInBuf[225]));
    AND2 select_163_Select_29_i1 (.O(n1_adj_1), .I0(state[7]), .I1(n5747));
    OR2 i3226 (.O(n6047), .I0(n6046), .I1(n6045));
    AND2 i2234 (.O(n5057), .I0(cnt[0]), .I1(cnt[1]));
    AND2 i3392 (.O(n6213), .I0(lcdRs_N_618), .I1(dataInBuf[224]));
    XOR2 i209 (.O(dispCount_5__N_347[3]), .I0(n3040), .I1(dispCount[3]));
    AND2 i3389 (.O(n6210), .I0(lcdRs_N_618), .I1(dataInBuf[222]));
    AND2 i3386 (.O(n6207), .I0(lcdRs_N_618), .I1(dataInBuf[221]));
    AND2 i3383 (.O(n6204), .I0(lcdRs_N_618), .I1(dataInBuf[220]));
    AND2 i3380 (.O(n6201), .I0(lcdRs_N_618), .I1(dataInBuf[219]));
    AND2 i3377 (.O(n6198), .I0(lcdRs_N_618), .I1(dataInBuf[218]));
    AND2 i3374 (.O(n6195), .I0(lcdRs_N_618), .I1(dataInBuf[217]));
    AND2 i3180 (.O(n6001), .I0(lcdRs_N_619), .I1(dataInBuf[150]));
    AND2 i3371 (.O(n6192), .I0(lcdRs_N_618), .I1(dataInBuf[216]));
    AND2 i3368 (.O(n6189), .I0(lcdRs_N_618), .I1(dataInBuf[214]));
    AND2 i3365 (.O(n6186), .I0(lcdRs_N_618), .I1(dataInBuf[213]));
    AND2 i3362 (.O(n6183), .I0(lcdRs_N_618), .I1(dataInBuf[212]));
    AND2 i3359 (.O(n6180), .I0(lcdRs_N_618), .I1(dataInBuf[211]));
    AND2 i3356 (.O(n6177), .I0(lcdRs_N_618), .I1(dataInBuf[210]));
    AND2 i3353 (.O(n6174), .I0(lcdRs_N_618), .I1(dataInBuf[209]));
    AND2 i3350 (.O(n6171), .I0(lcdRs_N_618), .I1(dataInBuf[208]));
    AND2 i3347 (.O(n6168), .I0(lcdRs_N_618), .I1(dataInBuf[206]));
    AND2 i3344 (.O(n6165), .I0(lcdRs_N_618), .I1(dataInBuf[205]));
    AND2 i3341 (.O(n6162), .I0(lcdRs_N_618), .I1(dataInBuf[204]));
    AND2 i3338 (.O(n6159), .I0(lcdRs_N_618), .I1(dataInBuf[203]));
    AND2 i3335 (.O(n6156), .I0(lcdRs_N_618), .I1(dataInBuf[202]));
    AND2 i3332 (.O(n6153), .I0(lcdRs_N_618), .I1(dataInBuf[201]));
    XOR2 i2343 (.O(n88), .I0(n5162), .I1(cnt[17]));
    AND2 i3329 (.O(n6150), .I0(lcdRs_N_618), .I1(dataInBuf[200]));
    AND2 i3326 (.O(n6147), .I0(lcdRs_N_618), .I1(dataInBuf[198]));
    AND2 i3323 (.O(n6144), .I0(lcdRs_N_618), .I1(dataInBuf[197]));
    AND2 i3320 (.O(n6141), .I0(lcdRs_N_618), .I1(dataInBuf[196]));
    AND2 i3317 (.O(n6138), .I0(lcdRs_N_618), .I1(dataInBuf[195]));
    AND2 i3314 (.O(n6135), .I0(lcdRs_N_618), .I1(dataInBuf[194]));
    AND2 i3311 (.O(n6132), .I0(lcdRs_N_618), .I1(dataInBuf[193]));
    OR2 i3181 (.O(n6002), .I0(n6001), .I1(n6000));
    AND2 i3308 (.O(n6129), .I0(lcdRs_N_618), .I1(dataInBuf[192]));
    AND2 i3305 (.O(n6126), .I0(lcdRs_N_618), .I1(dataInBuf[190]));
    AND2 i3302 (.O(n6123), .I0(lcdRs_N_618), .I1(dataInBuf[189]));
    AND2 i3299 (.O(n6120), .I0(lcdRs_N_618), .I1(dataInBuf[188]));
    AND2 i3296 (.O(n6117), .I0(lcdRs_N_618), .I1(dataInBuf[187]));
    AND2 i3293 (.O(n6114), .I0(lcdRs_N_618), .I1(dataInBuf[186]));
    AND2 i3290 (.O(n6111), .I0(lcdRs_N_618), .I1(dataInBuf[185]));
    AND2 i3183 (.O(n6004), .I0(lcdRs_N_619), .I1(dataInBuf[152]));
    AND2 i3287 (.O(n6108), .I0(lcdRs_N_618), .I1(dataInBuf[184]));
    AND2 i3284 (.O(n6105), .I0(lcdRs_N_618), .I1(dataInBuf[182]));
    AND2 i3281 (.O(n6102), .I0(lcdRs_N_618), .I1(dataInBuf[181]));
    AND2 i3278 (.O(n6099), .I0(lcdRs_N_618), .I1(dataInBuf[180]));
    AND2 i3275 (.O(n6096), .I0(lcdRs_N_618), .I1(dataInBuf[179]));
    AND2 i3272 (.O(n6093), .I0(lcdRs_N_618), .I1(dataInBuf[178]));
    AND2 i3269 (.O(n6090), .I0(lcdRs_N_618), .I1(dataInBuf[177]));
    AND2 i3266 (.O(n6087), .I0(lcdRs_N_618), .I1(dataInBuf[176]));
    AND2 i3263 (.O(n6084), .I0(lcdRs_N_618), .I1(dataInBuf[174]));
    AND2 i3260 (.O(n6081), .I0(lcdRs_N_618), .I1(dataInBuf[173]));
    AND2 i3257 (.O(n6078), .I0(lcdRs_N_618), .I1(dataInBuf[172]));
    AND2 i3254 (.O(n6075), .I0(lcdRs_N_618), .I1(dataInBuf[171]));
    AND2 i3251 (.O(n6072), .I0(lcdRs_N_618), .I1(dataInBuf[170]));
    AND2 i3248 (.O(n6069), .I0(lcdRs_N_618), .I1(dataInBuf[169]));
    AND2 i3245 (.O(n6066), .I0(lcdRs_N_618), .I1(dataInBuf[168]));
    AND2 i3242 (.O(n6063), .I0(lcdRs_N_618), .I1(dataInBuf[166]));
    AND2 i3239 (.O(n6060), .I0(lcdRs_N_618), .I1(dataInBuf[165]));
    AND2 i3236 (.O(n6057), .I0(lcdRs_N_618), .I1(dataInBuf[164]));
    AND2 i3233 (.O(n6054), .I0(lcdRs_N_618), .I1(dataInBuf[163]));
    AND2 i3230 (.O(n6051), .I0(lcdRs_N_618), .I1(dataInBuf[162]));
    AND2 i3227 (.O(n6048), .I0(lcdRs_N_618), .I1(dataInBuf[161]));
    OR2 i3184 (.O(n6005), .I0(n6004), .I1(n6003));
    AND2 i3224 (.O(n6045), .I0(lcdRs_N_618), .I1(dataInBuf[160]));
    AND2 i3221 (.O(n6042), .I0(lcdRs_N_618), .I1(dataInBuf[158]));
    AND2 i3218 (.O(n6039), .I0(lcdRs_N_618), .I1(dataInBuf[157]));
    AND2 i3215 (.O(n6036), .I0(lcdRs_N_618), .I1(dataInBuf[156]));
    AND2 i3212 (.O(n6033), .I0(lcdRs_N_618), .I1(dataInBuf[155]));
    AND2 i3209 (.O(n6030), .I0(lcdRs_N_618), .I1(dataInBuf[154]));
    AND2 i3206 (.O(n6027), .I0(lcdRs_N_618), .I1(dataInBuf[153]));
    AND2 i3203 (.O(n6024), .I0(lcdRs_N_618), .I1(dataInBuf[152]));
    AND2 i3200 (.O(n6021), .I0(lcdRs_N_618), .I1(dataInBuf[150]));
    AND2 i3197 (.O(n6018), .I0(lcdRs_N_618), .I1(dataInBuf[149]));
    AND2 i3194 (.O(n6015), .I0(lcdRs_N_618), .I1(dataInBuf[148]));
    AND2 i3191 (.O(n6012), .I0(lcdRs_N_618), .I1(dataInBuf[147]));
    AND2 i3188 (.O(n6009), .I0(lcdRs_N_618), .I1(dataInBuf[146]));
    AND2 i3185 (.O(n6006), .I0(lcdRs_N_618), .I1(dataInBuf[145]));
    AND2 i3182 (.O(n6003), .I0(lcdRs_N_618), .I1(dataInBuf[144]));
    AND2 i3179 (.O(n6000), .I0(lcdRs_N_618), .I1(dataInBuf[142]));
    AND2 i3176 (.O(n5997), .I0(lcdRs_N_618), .I1(dataInBuf[141]));
    AND2 i3173 (.O(n5994), .I0(lcdRs_N_618), .I1(dataInBuf[140]));
    AND2 i3170 (.O(n5991), .I0(lcdRs_N_618), .I1(dataInBuf[139]));
    AND2 i3167 (.O(n5988), .I0(lcdRs_N_618), .I1(dataInBuf[138]));
    AND2 i3164 (.O(n5985), .I0(lcdRs_N_618), .I1(dataInBuf[137]));
    OR2 i1537 (.O(lcdRs_N_617), .I0(lcdRs_N_620), .I1(lcdRs_N_618));
    AND2 i3161 (.O(n5982), .I0(lcdRs_N_618), .I1(dataInBuf[136]));
    AND2 i3158 (.O(n5979), .I0(lcdRs_N_618), .I1(dataInBuf[134]));
    AND2 i3155 (.O(n5976), .I0(lcdRs_N_618), .I1(dataInBuf[133]));
    AND2 i3152 (.O(n5973), .I0(lcdRs_N_618), .I1(dataInBuf[132]));
    AND2 i3149 (.O(n5970), .I0(lcdRs_N_618), .I1(dataInBuf[131]));
    AND2 i3146 (.O(n5967), .I0(lcdRs_N_618), .I1(dataInBuf[130]));
    AND2 i3143 (.O(n5964), .I0(lcdRs_N_618), .I1(dataInBuf[129]));
    AND2 i3186 (.O(n6007), .I0(lcdRs_N_619), .I1(dataInBuf[153]));
    AND2 i3140 (.O(n5961), .I0(lcdRs_N_618), .I1(dataInBuf[128]));
    AND2 i3137 (.O(n5958), .I0(lcdRs_N_618), .I1(dataInBuf[126]));
    AND2 i3294 (.O(n6115), .I0(lcdRs_N_619), .I1(dataInBuf[194]));
    OR2 select_163_Select_214_i9 (.O(n9_adj_380), .I0(n2_adj_379), .I1(n1_adj_378));
    AND2 select_163_Select_214_i2 (.O(n2_adj_379), .I0(state[6]), .I1(dataInBuf[206]));
    OR2 select_163_Select_218_i9 (.O(n9_adj_389), .I0(n2_adj_388), .I1(n1_adj_387));
    AND2 select_163_Select_217_i2 (.O(n2_adj_385), .I0(state[6]), .I1(dataInBuf[209]));
    AND2 i3134 (.O(n5955), .I0(lcdRs_N_618), .I1(dataInBuf[125]));
    AND2 select_163_Select_213_i2 (.O(n2_adj_377), .I0(state[6]), .I1(dataInBuf[205]));
    AND2 select_163_Select_156_i2 (.O(n2_adj_253), .I0(state[6]), .I1(dataInBuf[148]));
    AND2 i3131 (.O(n5952), .I0(lcdRs_N_618), .I1(dataInBuf[124]));
    OR2 i3295 (.O(n6116), .I0(n6115), .I1(n6114));
    AND2 i3128 (.O(n5949), .I0(lcdRs_N_618), .I1(dataInBuf[123]));
    OR2 i3418 (.O(n6239), .I0(n6238), .I1(n6237));
    OR2 select_163_Select_155_i9 (.O(n9_adj_251), .I0(n2_adj_250), .I1(n1_adj_249));
    AND2 i3036 (.O(n5857), .I0(lcdRs_N_619), .I1(dataInBuf[96]));
    AND2 i3125 (.O(n5946), .I0(lcdRs_N_618), .I1(dataInBuf[122]));
    AND2 i3420 (.O(n6241), .I0(lcdRs_N_619), .I1(dataInBuf[242]));
    AND2 select_163_Select_212_i2 (.O(n2_adj_375), .I0(state[6]), .I1(dataInBuf[204]));
    OR2 select_163_Select_211_i9 (.O(n9_adj_373), .I0(n2_adj_372), .I1(n1_adj_371));
    AND2 select_163_Select_218_i2 (.O(n2_adj_388), .I0(state[6]), .I1(dataInBuf[210]));
    AND2 i3122 (.O(n5943), .I0(lcdRs_N_618), .I1(dataInBuf[121]));
    OR2 i3421 (.O(n6242), .I0(n6241), .I1(n6240));
    AND2 select_163_Select_155_i2 (.O(n2_adj_250), .I0(state[6]), .I1(dataInBuf[147]));
    AND2 select_163_Select_211_i2 (.O(n2_adj_372), .I0(state[6]), .I1(dataInBuf[203]));
    OR2 select_163_Select_210_i9 (.O(n9_adj_370), .I0(n2_adj_369), .I1(n1_adj_368));
    AND2 select_163_Select_210_i2 (.O(n2_adj_369), .I0(state[6]), .I1(dataInBuf[202]));
    AND2 i3423 (.O(n6244), .I0(lcdRs_N_619), .I1(dataInBuf[243]));
    OR2 select_163_Select_209_i9 (.O(n9_adj_367), .I0(n2_adj_366), .I1(n1_adj_365));
    AND2 select_163_Select_209_i2 (.O(n2_adj_366), .I0(state[6]), .I1(dataInBuf[201]));
    AND2 select_163_Select_21_i1 (.O(n1_adj_11), .I0(state[7]), .I1(n5744));
    AND2 i3119 (.O(n5940), .I0(lcdRs_N_618), .I1(dataInBuf[120]));
    AND2 i3297 (.O(n6118), .I0(lcdRs_N_619), .I1(dataInBuf[195]));
    DFF cnt_171__i18 (.Q(cnt[18]), .D(n87), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i17 (.Q(cnt[17]), .D(n88), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i16 (.Q(cnt[16]), .D(n89), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i15 (.Q(cnt[15]), .D(n90), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i14 (.Q(cnt[14]), .D(n91), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i13 (.Q(cnt[13]), .D(n92), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i12 (.Q(cnt[12]), .D(n93), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i11 (.Q(cnt[11]), .D(n94), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i10 (.Q(cnt[10]), .D(n95), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i9 (.Q(cnt[9]), .D(n96), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i8 (.Q(cnt[8]), .D(n97), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i7 (.Q(cnt[7]), .D(n98), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i6 (.Q(cnt[6]), .D(n99), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i5 (.Q(cnt[5]), .D(n100), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i4 (.Q(cnt[4]), .D(n101), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i3 (.Q(cnt[3]), .D(n102), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i2 (.Q(cnt[2]), .D(n103), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFF cnt_171__i1 (.Q(cnt[1]), .D(n104), .CLK(clk_50m_c)) /* synthesis syn_use_carry_chain=1 */ ;   // lcd1602.v(43[24:31])
    DFFC dataInBuf_i0_i254 (.Q(dataInBuf[254]), .D(n9_adj_481), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i253 (.Q(dataInBuf[253]), .D(n5209), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i252 (.Q(dataInBuf[252]), .D(n9_adj_476), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i251 (.Q(dataInBuf[251]), .D(n9_adj_473), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i250 (.Q(dataInBuf[250]), .D(n9_adj_470), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i249 (.Q(dataInBuf[249]), .D(n9_adj_467), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i248 (.Q(dataInBuf[248]), .D(n9_adj_464), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i246 (.Q(dataInBuf[246]), .D(n9_adj_459), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3116 (.O(n5937), .I0(lcdRs_N_618), .I1(dataInBuf[118]));
    DFFC dataInBuf_i0_i245 (.Q(dataInBuf[245]), .D(n5659), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i244 (.Q(dataInBuf[244]), .D(n9_adj_454), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i243 (.Q(dataInBuf[243]), .D(n9_adj_451), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i242 (.Q(dataInBuf[242]), .D(n9_adj_448), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i241 (.Q(dataInBuf[241]), .D(n9_adj_445), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i240 (.Q(dataInBuf[240]), .D(n9_adj_442), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i238 (.Q(dataInBuf[238]), .D(n9_adj_439), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3113 (.O(n5934), .I0(lcdRs_N_618), .I1(dataInBuf[117]));
    DFFC dataInBuf_i0_i237 (.Q(dataInBuf[237]), .D(n5197), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i236 (.Q(dataInBuf[236]), .D(n9_adj_434), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i235 (.Q(dataInBuf[235]), .D(n9_adj_431), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i234 (.Q(dataInBuf[234]), .D(n9_adj_428), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i233 (.Q(dataInBuf[233]), .D(n9_adj_425), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i232 (.Q(dataInBuf[232]), .D(n9_adj_422), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i230 (.Q(dataInBuf[230]), .D(n9_adj_419), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i229 (.Q(dataInBuf[229]), .D(n5210), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i228 (.Q(dataInBuf[228]), .D(n9_adj_414), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i227 (.Q(dataInBuf[227]), .D(n9_adj_411), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i226 (.Q(dataInBuf[226]), .D(n9_adj_408), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i225 (.Q(dataInBuf[225]), .D(n9_adj_405), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i224 (.Q(dataInBuf[224]), .D(n9_adj_402), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i222 (.Q(dataInBuf[222]), .D(n9_adj_399), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i221 (.Q(dataInBuf[221]), .D(n5673), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i220 (.Q(dataInBuf[220]), .D(n5717), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i219 (.Q(dataInBuf[219]), .D(n9_adj_392), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i218 (.Q(dataInBuf[218]), .D(n9_adj_389), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i217 (.Q(dataInBuf[217]), .D(n9_adj_386), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i216 (.Q(dataInBuf[216]), .D(n9_adj_383), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i214 (.Q(dataInBuf[214]), .D(n9_adj_380), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i213 (.Q(dataInBuf[213]), .D(n5675), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i212 (.Q(dataInBuf[212]), .D(n5212), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i211 (.Q(dataInBuf[211]), .D(n9_adj_373), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i210 (.Q(dataInBuf[210]), .D(n9_adj_370), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i209 (.Q(dataInBuf[209]), .D(n9_adj_367), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i208 (.Q(dataInBuf[208]), .D(n5230), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i206 (.Q(dataInBuf[206]), .D(n9_adj_362), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3110 (.O(n5931), .I0(lcdRs_N_618), .I1(dataInBuf[116]));
    DFFC dataInBuf_i0_i205 (.Q(dataInBuf[205]), .D(n5715), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i204 (.Q(dataInBuf[204]), .D(n5677), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i203 (.Q(dataInBuf[203]), .D(n9_adj_355), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i202 (.Q(dataInBuf[202]), .D(n9_adj_352), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i201 (.Q(dataInBuf[201]), .D(n5214), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i200 (.Q(dataInBuf[200]), .D(n9_adj_347), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i198 (.Q(dataInBuf[198]), .D(n9_adj_344), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3107 (.O(n5928), .I0(lcdRs_N_618), .I1(dataInBuf[115]));
    DFFC dataInBuf_i0_i197 (.Q(dataInBuf[197]), .D(n5232), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i196 (.Q(dataInBuf[196]), .D(n5713), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i195 (.Q(dataInBuf[195]), .D(n9_adj_337), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i194 (.Q(dataInBuf[194]), .D(n9_adj_334), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i193 (.Q(dataInBuf[193]), .D(n5679), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i192 (.Q(dataInBuf[192]), .D(n5216), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i190 (.Q(dataInBuf[190]), .D(n9_adj_327), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i189 (.Q(dataInBuf[189]), .D(n5681), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i188 (.Q(dataInBuf[188]), .D(n5711), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i187 (.Q(dataInBuf[187]), .D(n9_adj_320), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i186 (.Q(dataInBuf[186]), .D(n5235), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i185 (.Q(dataInBuf[185]), .D(n9_adj_315), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i184 (.Q(dataInBuf[184]), .D(n9_adj_312), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i182 (.Q(dataInBuf[182]), .D(n9_adj_309), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i181 (.Q(dataInBuf[181]), .D(n5218), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i180 (.Q(dataInBuf[180]), .D(n5683), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3104 (.O(n5925), .I0(lcdRs_N_618), .I1(dataInBuf[114]));
    DFFC dataInBuf_i0_i179 (.Q(dataInBuf[179]), .D(n9_adj_302), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i178 (.Q(dataInBuf[178]), .D(n5709), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i177 (.Q(dataInBuf[177]), .D(n9_adj_297), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i176 (.Q(dataInBuf[176]), .D(n5237), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i174 (.Q(dataInBuf[174]), .D(n9_adj_292), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3101 (.O(n5922), .I0(lcdRs_N_618), .I1(dataInBuf[113]));
    DFFC dataInBuf_i0_i173 (.Q(dataInBuf[173]), .D(n5685), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i172 (.Q(dataInBuf[172]), .D(n5707), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i171 (.Q(dataInBuf[171]), .D(n9_adj_285), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3098 (.O(n5919), .I0(lcdRs_N_618), .I1(dataInBuf[112]));
    DFFC dataInBuf_i0_i170 (.Q(dataInBuf[170]), .D(n5239), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i169 (.Q(dataInBuf[169]), .D(n5221), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i168 (.Q(dataInBuf[168]), .D(n9_adj_278), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i166 (.Q(dataInBuf[166]), .D(n9_adj_275), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3095 (.O(n5916), .I0(lcdRs_N_618), .I1(dataInBuf[110]));
    DFFC dataInBuf_i0_i165 (.Q(dataInBuf[165]), .D(n5687), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i164 (.Q(dataInBuf[164]), .D(n5222), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i163 (.Q(dataInBuf[163]), .D(n9_adj_268), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i162 (.Q(dataInBuf[162]), .D(n5689), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i161 (.Q(dataInBuf[161]), .D(n5223), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i160 (.Q(dataInBuf[160]), .D(n5242), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i158 (.Q(dataInBuf[158]), .D(n9_adj_259), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i157 (.Q(dataInBuf[157]), .D(n5224), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i156 (.Q(dataInBuf[156]), .D(n9_adj_254), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i155 (.Q(dataInBuf[155]), .D(n9_adj_251), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i154 (.Q(dataInBuf[154]), .D(n9_adj_248), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i153 (.Q(dataInBuf[153]), .D(n9_adj_245), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i152 (.Q(dataInBuf[152]), .D(n9_adj_242), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i150 (.Q(dataInBuf[150]), .D(n9_adj_239), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i149 (.Q(dataInBuf[149]), .D(n5691), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i148 (.Q(dataInBuf[148]), .D(n9_adj_234), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i147 (.Q(dataInBuf[147]), .D(n9_adj_231), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i146 (.Q(dataInBuf[146]), .D(n9_adj_228), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i145 (.Q(dataInBuf[145]), .D(n9_adj_225), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i144 (.Q(dataInBuf[144]), .D(n9_adj_222), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i142 (.Q(dataInBuf[142]), .D(n9_adj_219), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i141 (.Q(dataInBuf[141]), .D(n5196), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i140 (.Q(dataInBuf[140]), .D(n9_adj_214), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i139 (.Q(dataInBuf[139]), .D(n9_adj_211), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i138 (.Q(dataInBuf[138]), .D(n9_adj_208), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i137 (.Q(dataInBuf[137]), .D(n9_adj_205), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i136 (.Q(dataInBuf[136]), .D(n9_adj_202), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i134 (.Q(dataInBuf[134]), .D(n9_adj_199), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3092 (.O(n5913), .I0(lcdRs_N_618), .I1(dataInBuf[109]));
    DFFC dataInBuf_i0_i133 (.Q(dataInBuf[133]), .D(n5244), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i132 (.Q(dataInBuf[132]), .D(n9_adj_194), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i131 (.Q(dataInBuf[131]), .D(n9_adj_191), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i130 (.Q(dataInBuf[130]), .D(n9_adj_188), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i129 (.Q(dataInBuf[129]), .D(n9_adj_185), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i128 (.Q(dataInBuf[128]), .D(n9_adj_182), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i126 (.Q(dataInBuf[126]), .D(n9_adj_179), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3089 (.O(n5910), .I0(lcdRs_N_618), .I1(dataInBuf[108]));
    DFFC dataInBuf_i0_i125 (.Q(dataInBuf[125]), .D(n5693), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i124 (.Q(dataInBuf[124]), .D(n9_adj_174), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i123 (.Q(dataInBuf[123]), .D(n9_adj_171), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i122 (.Q(dataInBuf[122]), .D(n9_adj_168), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i121 (.Q(dataInBuf[121]), .D(n9_adj_165), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i120 (.Q(dataInBuf[120]), .D(n9_adj_162), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i118 (.Q(dataInBuf[118]), .D(n9_adj_159), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3086 (.O(n5907), .I0(lcdRs_N_618), .I1(dataInBuf[107]));
    DFFC dataInBuf_i0_i117 (.Q(dataInBuf[117]), .D(n5671), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i116 (.Q(dataInBuf[116]), .D(n9_adj_154), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i115 (.Q(dataInBuf[115]), .D(n9_adj_151), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i114 (.Q(dataInBuf[114]), .D(n9_adj_148), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i113 (.Q(dataInBuf[113]), .D(n9_adj_145), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i112 (.Q(dataInBuf[112]), .D(n9_adj_142), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i110 (.Q(dataInBuf[110]), .D(n9_adj_139), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i109 (.Q(dataInBuf[109]), .D(n5246), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i108 (.Q(dataInBuf[108]), .D(n9_adj_134), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i107 (.Q(dataInBuf[107]), .D(n9_adj_131), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i106 (.Q(dataInBuf[106]), .D(n9_adj_128), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i105 (.Q(dataInBuf[105]), .D(n9_adj_125), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i104 (.Q(dataInBuf[104]), .D(n9_adj_122), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i102 (.Q(dataInBuf[102]), .D(n9_adj_119), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i101 (.Q(dataInBuf[101]), .D(n5199), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i100 (.Q(dataInBuf[100]), .D(n9_adj_114), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i99 (.Q(dataInBuf[99]), .D(n9_adj_111), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i98 (.Q(dataInBuf[98]), .D(n9_adj_108), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i97 (.Q(dataInBuf[97]), .D(n9_adj_105), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i96 (.Q(dataInBuf[96]), .D(n9_adj_102), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i94 (.Q(dataInBuf[94]), .D(n9_adj_99), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3083 (.O(n5904), .I0(lcdRs_N_618), .I1(dataInBuf[106]));
    DFFC dataInBuf_i0_i93 (.Q(dataInBuf[93]), .D(n5695), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i92 (.Q(dataInBuf[92]), .D(n5669), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i91 (.Q(dataInBuf[91]), .D(n5248), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i90 (.Q(dataInBuf[90]), .D(n9_adj_90), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i89 (.Q(dataInBuf[89]), .D(n9_adj_87), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i88 (.Q(dataInBuf[88]), .D(n9_adj_84), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i86 (.Q(dataInBuf[86]), .D(n9_adj_81), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i85 (.Q(dataInBuf[85]), .D(n5201), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3080 (.O(n5901), .I0(lcdRs_N_618), .I1(dataInBuf[105]));
    DFFC dataInBuf_i0_i84 (.Q(dataInBuf[84]), .D(n3753), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i83 (.Q(dataInBuf[83]), .D(n4), .CLK(ledEN_c), .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i82 (.Q(dataInBuf[82]), .D(n9_adj_76), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i81 (.Q(dataInBuf[81]), .D(n9_adj_73), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i80 (.Q(dataInBuf[80]), .D(n5697), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i78 (.Q(dataInBuf[78]), .D(n5667), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3077 (.O(n5898), .I0(lcdRs_N_618), .I1(dataInBuf[104]));
    DFFC dataInBuf_i0_i77 (.Q(dataInBuf[77]), .D(n9_adj_66), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i74 (.Q(dataInBuf[74]), .D(n9_adj_63), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i73 (.Q(dataInBuf[73]), .D(n9_adj_60), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i72 (.Q(dataInBuf[72]), .D(n5250), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i70 (.Q(dataInBuf[70]), .D(n5203), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3074 (.O(n5895), .I0(lcdRs_N_618), .I1(dataInBuf[102]));
    DFFC dataInBuf_i0_i69 (.Q(dataInBuf[69]), .D(n9_adj_53), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i66 (.Q(dataInBuf[66]), .D(n9_adj_50), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3071 (.O(n5892), .I0(lcdRs_N_618), .I1(dataInBuf[101]));
    DFFC dataInBuf_i0_i65 (.Q(dataInBuf[65]), .D(n5699), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i64 (.Q(dataInBuf[64]), .D(n9_adj_45), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i62 (.Q(dataInBuf[62]), .D(n5665), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i61 (.Q(dataInBuf[61]), .D(n9_adj_40), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i58 (.Q(dataInBuf[58]), .D(n9_adj_37), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3068 (.O(n5889), .I0(lcdRs_N_618), .I1(dataInBuf[100]));
    AND2 i3065 (.O(n5886), .I0(lcdRs_N_618), .I1(dataInBuf[99]));
    DFFC dataInBuf_i0_i57 (.Q(dataInBuf[57]), .D(n5701), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i56 (.Q(dataInBuf[56]), .D(n5205), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i54 (.Q(dataInBuf[54]), .D(n5253), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i53 (.Q(dataInBuf[53]), .D(n9_adj_28), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i50 (.Q(dataInBuf[50]), .D(n5255), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3062 (.O(n5883), .I0(lcdRs_N_618), .I1(dataInBuf[98]));
    DFFC dataInBuf_i0_i49 (.Q(dataInBuf[49]), .D(n9_adj_14), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i48 (.Q(dataInBuf[48]), .D(n3739), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i46 (.Q(dataInBuf[46]), .D(n5663), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3059 (.O(n5880), .I0(lcdRs_N_618), .I1(dataInBuf[97]));
    DFFC dataInBuf_i0_i45 (.Q(dataInBuf[45]), .D(n9_adj_24), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i42 (.Q(dataInBuf[42]), .D(n5207), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i41 (.Q(dataInBuf[41]), .D(n9), .CLK(ledEN_c), .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i38 (.Q(dataInBuf[38]), .D(n4_adj_461), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i37 (.Q(dataInBuf[37]), .D(n9_adj_17), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i34 (.Q(dataInBuf[34]), .D(n3733), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i33 (.Q(dataInBuf[33]), .D(n4_adj_460), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i29 (.Q(dataInBuf[29]), .D(n5259), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    DFFC dataInBuf_i0_i21 (.Q(dataInBuf[21]), .D(n5661), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3056 (.O(n5877), .I0(lcdRs_N_618), .I1(dataInBuf[96]));
    AND2 i3053 (.O(n5874), .I0(lcdRs_N_618), .I1(dataInBuf[94]));
    DFFC dataInBuf_i0_i13 (.Q(dataInBuf[13]), .D(n5703), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3050 (.O(n5871), .I0(lcdRs_N_618), .I1(dataInBuf[93]));
    AND2 i3047 (.O(n5868), .I0(lcdRs_N_618), .I1(dataInBuf[92]));
    AND2 i3044 (.O(n5865), .I0(lcdRs_N_618), .I1(dataInBuf[91]));
    AND2 i3041 (.O(n5862), .I0(lcdRs_N_618), .I1(dataInBuf[90]));
    DFFC dataInBuf_i0_i5 (.Q(dataInBuf[5]), .D(n3000), .CLK(ledEN_c), 
         .CE(n3805));   // lcd1602.v(62[14] 139[12])
    AND2 i3038 (.O(n5859), .I0(lcdRs_N_618), .I1(dataInBuf[89]));
    OR2 i3187 (.O(n6008), .I0(n6007), .I1(n6006));
    AND2 i3035 (.O(n5856), .I0(lcdRs_N_618), .I1(dataInBuf[88]));
    AND2 i3032 (.O(n5853), .I0(lcdRs_N_618), .I1(dataInBuf[86]));
    DFFS state_FSM_i7 (.Q(state[0]), .D(n2212), .CLK(ledEN_c), .S(reset_c));   // lcd1602.v(63[13] 138[20])
    AND2 i3029 (.O(n5850), .I0(lcdRs_N_618), .I1(dataInBuf[85]));
    OR3 i1_adj_29 (.O(n5665), .I0(n1_adj_41), .I1(n2_adj_42), .I2(state[0]));
    AND2 select_163_Select_208_i2 (.O(n2_adj_364), .I0(state[6]), .I1(dataInBuf[200]));
    OR2 i3298 (.O(n6119), .I0(n6118), .I1(n6117));
    OR2 i2956 (.O(n5777), .I0(n5776), .I1(n5775));
    AND2 i3300 (.O(n6121), .I0(lcdRs_N_619), .I1(dataInBuf[196]));
    OR2 i3301 (.O(n6122), .I0(n6121), .I1(n6120));
    AND2 i2958 (.O(n5779), .I0(lcdRs_N_619), .I1(dataInBuf[57]));
    AND2 i3303 (.O(n6124), .I0(lcdRs_N_619), .I1(dataInBuf[197]));
    OR2 i3304 (.O(n6125), .I0(n6124), .I1(n6123));
    OR2 select_163_Select_206_i9 (.O(n9_adj_362), .I0(n2_adj_361), .I1(n1_adj_360));
    OR2 i2959 (.O(n5780), .I0(n5779), .I1(n5778));
    AND2 i3306 (.O(n6127), .I0(lcdRs_N_619), .I1(dataInBuf[198]));
    OR2 i3307 (.O(n6128), .I0(n6127), .I1(n6126));
    AND2 select_163_Select_206_i2 (.O(n2_adj_361), .I0(state[6]), .I1(dataInBuf[198]));
    AND2 i2961 (.O(n5782), .I0(lcdRs_N_619), .I1(dataInBuf[58]));
    AND2 i3309 (.O(n6130), .I0(lcdRs_N_619), .I1(dataInBuf[200]));
    OR2 i2962 (.O(n5783), .I0(n5782), .I1(n5781));
    OR2 i3310 (.O(n6131), .I0(n6130), .I1(n6129));
    AND2 i3312 (.O(n6133), .I0(lcdRs_N_619), .I1(dataInBuf[201]));
    XOR2 i2350 (.O(n87), .I0(n5169), .I1(cnt[18]));
    AND2 select_163_Select_205_i2 (.O(n2_adj_359), .I0(state[6]), .I1(dataInBuf[197]));
    XOR2 i2252 (.O(n101), .I0(n5071), .I1(cnt[4]));
    AND2 i2346 (.O(n5169), .I0(n5162), .I1(cnt[17]));
    OR3 i2_adj_30 (.O(n5257), .I0(state[6]), .I1(n5650), .I2(state[4]));
    AND2 i2262 (.O(n5085), .I0(n5078), .I1(cnt[5]));
    AND2 i2964 (.O(n5785), .I0(lcdRs_N_619), .I1(dataInBuf[61]));
    XOR2 i2357 (.O(n86), .I0(n5176), .I1(cnt[19]));
    OR3 i1_adj_31 (.O(n5701), .I0(n2_adj_34), .I1(n1_adj_33), .I2(state[0]));
    AND2 select_163_Select_204_i2 (.O(n2_adj_357), .I0(state[6]), .I1(dataInBuf[196]));
    OR2 i3313 (.O(n6134), .I0(n6133), .I1(n6132));
    AND2 i3315 (.O(n6136), .I0(lcdRs_N_619), .I1(dataInBuf[202]));
    OR2 select_163_Select_203_i9 (.O(n9_adj_355), .I0(n2_adj_354), .I1(n1_adj_353));
    OR2 i2965 (.O(n5786), .I0(n5785), .I1(n5784));
    AND2 select_163_Select_203_i2 (.O(n2_adj_354), .I0(state[6]), .I1(dataInBuf[195]));
    OR2 select_163_Select_202_i9 (.O(n9_adj_352), .I0(n2_adj_351), .I1(n1_adj_350));
    OR3 i2_adj_32 (.O(n5209), .I0(n1_adj_477), .I1(n2_adj_478), .I2(state[0]));
    AND2 i2967 (.O(n5788), .I0(lcdRs_N_619), .I1(dataInBuf[62]));
    AND2 select_163_Select_202_i2 (.O(n2_adj_351), .I0(state[6]), .I1(dataInBuf[194]));
    OR2 i2968 (.O(n5789), .I0(n5788), .I1(n5787));
    OR2 i3316 (.O(n6137), .I0(n6136), .I1(n6135));
    AND2 i2970 (.O(n5791), .I0(lcdRs_N_619), .I1(dataInBuf[64]));
    AND2 select_163_Select_201_i2 (.O(n2_adj_349), .I0(state[6]), .I1(dataInBuf[193]));
    AND2 i3318 (.O(n6139), .I0(lcdRs_N_619), .I1(dataInBuf[203]));
    OR2 select_163_Select_200_i9 (.O(n9_adj_347), .I0(n2_adj_346), .I1(n1_adj_345));
    OR2 i3319 (.O(n6140), .I0(n6139), .I1(n6138));
    AND2 select_163_Select_200_i2 (.O(n2_adj_346), .I0(state[6]), .I1(dataInBuf[192]));
    OR2 i2971 (.O(n5792), .I0(n5791), .I1(n5790));
    AND2 i3026 (.O(n5847), .I0(lcdRs_N_618), .I1(dataInBuf[84]));
    AND2 i3321 (.O(n6142), .I0(lcdRs_N_619), .I1(dataInBuf[204]));
    OR2 i3322 (.O(n6143), .I0(n6142), .I1(n6141));
    OR2 select_163_Select_198_i9 (.O(n9_adj_344), .I0(n2_adj_343), .I1(n1_adj_342));
    AND2 i2973 (.O(n5794), .I0(lcdRs_N_619), .I1(dataInBuf[65]));
    AND2 select_163_Select_198_i2 (.O(n2_adj_343), .I0(state[6]), .I1(dataInBuf[190]));
    OR3 i2_adj_33 (.O(n5207), .I0(n1_adj_2), .I1(n2_adj_3), .I2(state[0]));
    AND2 select_163_Select_197_i2 (.O(n2_adj_341), .I0(state[6]), .I1(dataInBuf[189]));
    AND2 i3324 (.O(n6145), .I0(lcdRs_N_619), .I1(dataInBuf[205]));
    OR2 i3325 (.O(n6146), .I0(n6145), .I1(n6144));
    OR2 i2974 (.O(n5795), .I0(n5794), .I1(n5793));
    AND2 select_163_Select_196_i2 (.O(n2_adj_339), .I0(state[6]), .I1(dataInBuf[188]));
    OR2 select_163_Select_195_i9 (.O(n9_adj_337), .I0(n2_adj_336), .I1(n1_adj_335));
    AND2 select_163_Select_195_i2 (.O(n2_adj_336), .I0(state[6]), .I1(dataInBuf[187]));
    OR2 select_163_Select_194_i9 (.O(n9_adj_334), .I0(n2_adj_333), .I1(n1_adj_332));
    AND2 select_163_Select_194_i2 (.O(n2_adj_333), .I0(state[6]), .I1(dataInBuf[186]));
    AND2 i2976 (.O(n5797), .I0(lcdRs_N_619), .I1(dataInBuf[66]));
    OR3 i2_adj_34 (.O(n5205), .I0(n1_adj_31), .I1(n2_adj_32), .I2(state[0]));
    AND2 select_163_Select_193_i2 (.O(n2_adj_331), .I0(state[6]), .I1(dataInBuf[185]));
    AND2 i3327 (.O(n6148), .I0(lcdRs_N_619), .I1(dataInBuf[206]));
    OR2 i3328 (.O(n6149), .I0(n6148), .I1(n6147));
    OR2 i2977 (.O(n5798), .I0(n5797), .I1(n5796));
    AND2 i1592 (.O(n2159), .I0(n2185), .I1(dispCount_5__N_347[0]));
    AND2 select_163_Select_192_i2 (.O(n2_adj_329), .I0(state[6]), .I1(dataInBuf[184]));
    AND2 i2979 (.O(n5800), .I0(lcdRs_N_619), .I1(dataInBuf[69]));
    AND2 i3330 (.O(n6151), .I0(lcdRs_N_619), .I1(dataInBuf[208]));
    OR2 select_163_Select_190_i9 (.O(n9_adj_327), .I0(n2_adj_326), .I1(n1_adj_325));
    AND2 select_163_Select_190_i2 (.O(n2_adj_326), .I0(state[6]), .I1(dataInBuf[182]));
    AND2 select_163_Select_189_i2 (.O(n2_adj_324), .I0(state[6]), .I1(dataInBuf[181]));
    OR2 i3331 (.O(n6152), .I0(n6151), .I1(n6150));
    OR2 i2980 (.O(n5801), .I0(n5800), .I1(n5799));
    AND2 select_163_Select_188_i2 (.O(n2_adj_322), .I0(state[6]), .I1(dataInBuf[180]));
    AND2 i3333 (.O(n6154), .I0(lcdRs_N_619), .I1(dataInBuf[209]));
    OR2 select_163_Select_187_i9 (.O(n9_adj_320), .I0(n2_adj_319), .I1(n1_adj_318));
    AND2 select_163_Select_187_i2 (.O(n2_adj_319), .I0(state[6]), .I1(dataInBuf[179]));
    OR2 i3334 (.O(n6155), .I0(n6154), .I1(n6153));
    OR3 i2_adj_35 (.O(n5203), .I0(n1_adj_54), .I1(n2_adj_55), .I2(state[0]));
    AND2 select_163_Select_186_i2 (.O(n2_adj_317), .I0(state[6]), .I1(dataInBuf[178]));
    OR2 select_163_Select_185_i9 (.O(n9_adj_315), .I0(n2_adj_314), .I1(n1_adj_313));
    AND2 i3336 (.O(n6157), .I0(lcdRs_N_619), .I1(dataInBuf[210]));
    AND2 select_163_Select_185_i2 (.O(n2_adj_314), .I0(state[6]), .I1(dataInBuf[177]));
    OR2 select_163_Select_184_i9 (.O(n9_adj_312), .I0(n2_adj_311), .I1(n1_adj_310));
    AND2 i2353 (.O(n5176), .I0(n5169), .I1(cnt[18]));
    AND2 select_163_Select_184_i2 (.O(n2_adj_311), .I0(state[6]), .I1(dataInBuf[176]));
    AND2 i2269 (.O(n5092), .I0(n5085), .I1(cnt[6]));
    AND2 i2982 (.O(n5803), .I0(lcdRs_N_619), .I1(dataInBuf[70]));
    OR2 i3337 (.O(n6158), .I0(n6157), .I1(n6156));
    OR2 select_163_Select_182_i9 (.O(n9_adj_309), .I0(n2_adj_308), .I1(n1_adj_307));
    AND2 select_163_Select_182_i2 (.O(n2_adj_308), .I0(state[6]), .I1(dataInBuf[174]));
    OR2 i2983 (.O(n5804), .I0(n5803), .I1(n5802));
    AND2 i3339 (.O(n6160), .I0(lcdRs_N_619), .I1(dataInBuf[211]));
    AND2 i2985 (.O(n5806), .I0(lcdRs_N_619), .I1(dataInBuf[72]));
    AND2 select_163_Select_181_i2 (.O(n2_adj_306), .I0(state[6]), .I1(dataInBuf[173]));
    OR2 i3340 (.O(n6161), .I0(n6160), .I1(n6159));
    AND2 select_163_Select_180_i2 (.O(n2_adj_304), .I0(state[6]), .I1(dataInBuf[172]));
    OR2 select_163_Select_179_i9 (.O(n9_adj_302), .I0(n2_adj_301), .I1(n1_adj_300));
    AND2 i3342 (.O(n6163), .I0(lcdRs_N_619), .I1(dataInBuf[212]));
    AND2 select_163_Select_179_i2 (.O(n2_adj_301), .I0(state[6]), .I1(dataInBuf[171]));
    AND2 i3471 (.O(n6292), .I0(n6285), .I1(n20));
    AND2 i3468 (.O(n6289), .I0(n6285), .I1(n44));
    OR2 i3343 (.O(n6164), .I0(n6163), .I1(n6162));
    AND2 i3345 (.O(n6166), .I0(lcdRs_N_619), .I1(dataInBuf[213]));
    AND2 select_163_Select_178_i2 (.O(n2_adj_299), .I0(state[6]), .I1(dataInBuf[170]));
    OR2 select_163_Select_177_i9 (.O(n9_adj_297), .I0(n2_adj_296), .I1(n1_adj_295));
    OR3 i2_adj_36 (.O(n5201), .I0(n1_adj_77), .I1(n2_adj_78), .I2(state[0]));
    OR2 i2986 (.O(n5807), .I0(n5806), .I1(n5805));
    AND2 select_163_Select_177_i2 (.O(n2_adj_296), .I0(state[6]), .I1(dataInBuf[169]));
    AND2 i1570 (.O(n44), .I0(state[2]), .I1(n14_adj_6));
    AND2 i1_adj_37 (.O(n3731), .I0(n16), .I1(n3729));
    AND2 i2988 (.O(n5809), .I0(lcdRs_N_619), .I1(dataInBuf[73]));
    AND2 select_163_Select_176_i2 (.O(n2_adj_294), .I0(state[6]), .I1(dataInBuf[168]));
    OR2 i3346 (.O(n6167), .I0(n6166), .I1(n6165));
    OR2 i1568 (.O(n33), .I0(n4374), .I1(dataInBuf[254]));
    AND2 i3348 (.O(n6169), .I0(lcdRs_N_619), .I1(dataInBuf[214]));
    OR2 i2989 (.O(n5810), .I0(n5809), .I1(n5808));
    OR2 select_163_Select_174_i9 (.O(n9_adj_292), .I0(n2_adj_291), .I1(n1_adj_290));
    OR2 i1562 (.O(n3637), .I0(n3012), .I1(n5719));
    AND2 i1561 (.O(n2199), .I0(n40), .I1(n33));
    OR3 i2_adj_38 (.O(n5199), .I0(n1_adj_115), .I1(n2_adj_116), .I2(state[0]));
    OR2 i1560 (.O(n3117), .I0(state[4]), .I1(state[3]));
    AND2 select_163_Select_174_i2 (.O(n2_adj_291), .I0(state[6]), .I1(dataInBuf[166]));
    AND2 i2991 (.O(n5812), .I0(lcdRs_N_619), .I1(dataInBuf[74]));
    AND2 i3023 (.O(n5844), .I0(lcdRs_N_618), .I1(dataInBuf[83]));
    AND2 i1559 (.O(n2160), .I0(n2185), .I1(dispCount_5__N_347[1]));
    AND2 i1558 (.O(n2161), .I0(n2185), .I1(dispCount_5__N_347[2]));
    AND2 i1557 (.O(n2162), .I0(n2185), .I1(dispCount_5__N_347[3]));
    OR3 i1_adj_39 (.O(n5703), .I0(n2_adj_19), .I1(n1_adj_18), .I2(state[0]));
    AND2 i1556 (.O(n2163), .I0(n2185), .I1(dispCount_5__N_347[4]));
    OR2 i3349 (.O(n6170), .I0(n6169), .I1(n6168));
    XOR2 i1_adj_40 (.O(ledEN_N_622), .I0(n5194), .I1(ledEN_c));
    AND2 select_163_Select_173_i2 (.O(n2_adj_289), .I0(state[6]), .I1(dataInBuf[165]));
    AND2 i3351 (.O(n6172), .I0(lcdRs_N_619), .I1(dataInBuf[216]));
    AND2 i3020 (.O(n5841), .I0(lcdRs_N_618), .I1(dataInBuf[82]));
    OR3 i2_adj_41 (.O(n5197), .I0(n1_adj_435), .I1(n2_adj_436), .I2(state[0]));
    AND2 i2919 (.O(n5740), .I0(lcdRs_N_619), .I1(dataInBuf[13]));
    OR2 i3352 (.O(n6173), .I0(n6172), .I1(n6171));
    AND2 i3354 (.O(n6175), .I0(lcdRs_N_619), .I1(dataInBuf[217]));
    OR2 i3355 (.O(n6176), .I0(n6175), .I1(n6174));
    OR2 i1_adj_42 (.O(n3739), .I0(n5726), .I1(state[0]));
    OR3 i1_adj_43 (.O(n5667), .I0(n1_adj_67), .I1(n2_adj_68), .I2(state[0]));
    AND2 select_163_Select_172_i2 (.O(n2_adj_287), .I0(state[6]), .I1(dataInBuf[164]));
    AND2 i2922 (.O(n5743), .I0(lcdRs_N_619), .I1(dataInBuf[21]));
    OR2 i2992 (.O(n5813), .I0(n5812), .I1(n5811));
    AND2 i3017 (.O(n5838), .I0(lcdRs_N_618), .I1(dataInBuf[81]));
    OR2 select_163_Select_171_i9 (.O(n9_adj_285), .I0(n2_adj_284), .I1(n1_adj_283));
    AND2 i2994 (.O(n5815), .I0(lcdRs_N_619), .I1(dataInBuf[77]));
    OR2 i2995 (.O(n5816), .I0(n5815), .I1(n5814));
    AND2 i3357 (.O(n6178), .I0(lcdRs_N_619), .I1(dataInBuf[218]));
    AND2 select_163_Select_171_i2 (.O(n2_adj_284), .I0(state[6]), .I1(dataInBuf[163]));
    AND2 i2997 (.O(n5818), .I0(lcdRs_N_619), .I1(dataInBuf[78]));
    AND2 i2311 (.O(n5134), .I0(n5127), .I1(cnt[12]));
    OR4 i3_adj_44 (.O(n3800), .I0(dispCount[1]), .I1(dispCount[2]), .I2(dispCount[0]), 
        .I3(dispCount[3]));
    OR2 i3358 (.O(n6179), .I0(n6178), .I1(n6177));
    OR2 i2998 (.O(n5819), .I0(n5818), .I1(n5817));
    OR3 i1_adj_45 (.O(n5707), .I0(n1_adj_286), .I1(n2_adj_287), .I2(state[0]));
    AND2 i3360 (.O(n6181), .I0(lcdRs_N_619), .I1(dataInBuf[219]));
    AND2 select_163_Select_170_i2 (.O(n2_adj_282), .I0(state[6]), .I1(dataInBuf[162]));
    AND2 i3000 (.O(n5821), .I0(lcdRs_N_619), .I1(dataInBuf[80]));
    OR2 i3361 (.O(n6182), .I0(n6181), .I1(n6180));
    AND2 i3363 (.O(n6184), .I0(lcdRs_N_619), .I1(dataInBuf[220]));
    OR2 i1_adj_46 (.O(n3753), .I0(n5728), .I1(state[0]));
    OR2 i3364 (.O(n6185), .I0(n6184), .I1(n6183));
    AND4 i3_adj_47 (.O(n3012), .I0(n3729), .I1(n1_adj_10), .I2(state[7]), 
         .I3(dispCount[4]));
    AND2 select_163_Select_169_i2 (.O(n2_adj_280), .I0(state[6]), .I1(dataInBuf[161]));
    OR2 i3001 (.O(n5822), .I0(n5821), .I1(n5820));
    AND2 i3366 (.O(n6187), .I0(lcdRs_N_619), .I1(dataInBuf[221]));
    OR2 i3367 (.O(n6188), .I0(n6187), .I1(n6186));
    OR3 i1_adj_48 (.O(n5709), .I0(n1_adj_298), .I1(n2_adj_299), .I2(state[0]));
    OR2 select_163_Select_168_i9 (.O(n9_adj_278), .I0(n2_adj_277), .I1(n1_adj_276));
    OR3 i2_adj_49 (.O(n5224), .I0(n1_adj_255), .I1(n2_adj_256), .I2(state[0]));
    AND2 i3369 (.O(n6190), .I0(lcdRs_N_619), .I1(dataInBuf[222]));
    AND2 select_163_Select_168_i2 (.O(n2_adj_277), .I0(state[6]), .I1(dataInBuf[160]));
    AND2 i3003 (.O(n5824), .I0(lcdRs_N_619), .I1(dataInBuf[81]));
    OR2 i3004 (.O(n5825), .I0(n5824), .I1(n5823));
    OR2 i3370 (.O(n6191), .I0(n6190), .I1(n6189));
    AND2 i3372 (.O(n6193), .I0(lcdRs_N_619), .I1(dataInBuf[224]));
    OR3 i2_adj_50 (.O(n5230), .I0(n1_adj_363), .I1(state[0]), .I2(n2_adj_364));
    AND2 i3006 (.O(n5827), .I0(lcdRs_N_619), .I1(dataInBuf[82]));
    OR2 i3373 (.O(n6194), .I0(n6193), .I1(n6192));
    OR2 i3007 (.O(n5828), .I0(n5827), .I1(n5826));
    AND2 i3375 (.O(n6196), .I0(lcdRs_N_619), .I1(dataInBuf[225]));
    OR3 i2_adj_51 (.O(n5232), .I0(n1_adj_340), .I1(state[0]), .I2(n2_adj_341));
    OR2 select_163_Select_166_i9 (.O(n9_adj_275), .I0(n2_adj_274), .I1(n1_adj_273));
    OR2 i3376 (.O(n6197), .I0(n6196), .I1(n6195));
    AND2 i3378 (.O(n6199), .I0(lcdRs_N_619), .I1(dataInBuf[226]));
    AND2 select_163_Select_166_i2 (.O(n2_adj_274), .I0(state[6]), .I1(dataInBuf[158]));
    OR2 i3379 (.O(n6200), .I0(n6199), .I1(n6198));
    AND2 i3009 (.O(n5830), .I0(lcdRs_N_619), .I1(dataInBuf[85]));
    OR3 i2_adj_52 (.O(n5223), .I0(n1_adj_262), .I1(n2_adj_263), .I2(state[0]));
    AND2 i3381 (.O(n6202), .I0(lcdRs_N_619), .I1(dataInBuf[227]));
    OR3 i1_adj_53 (.O(n5711), .I0(n1_adj_321), .I1(n2_adj_322), .I2(state[0]));
    OR3 i2_adj_54 (.O(n5235), .I0(n1_adj_316), .I1(state[0]), .I2(n2_adj_317));
    OR2 i3010 (.O(n5831), .I0(n5830), .I1(n5829));
    OR2 i3382 (.O(n6203), .I0(n6202), .I1(n6201));
    AND2 select_163_Select_165_i2 (.O(n2_adj_272), .I0(state[6]), .I1(dataInBuf[157]));
    AND2 i3012 (.O(n5833), .I0(lcdRs_N_619), .I1(dataInBuf[86]));
    OR2 i3013 (.O(n5834), .I0(n5833), .I1(n5832));
    AND2 i3384 (.O(n6205), .I0(lcdRs_N_619), .I1(dataInBuf[228]));
    OR3 i2_adj_55 (.O(n5237), .I0(n1_adj_293), .I1(state[0]), .I2(n2_adj_294));
    AND2 i3015 (.O(n5836), .I0(lcdRs_N_619), .I1(dataInBuf[88]));
    OR2 i3385 (.O(n6206), .I0(n6205), .I1(n6204));
    AND2 select_163_Select_164_i2 (.O(n2_adj_270), .I0(state[6]), .I1(dataInBuf[156]));
    OR2 i3016 (.O(n5837), .I0(n5836), .I1(n5835));
    AND2 i3387 (.O(n6208), .I0(lcdRs_N_619), .I1(dataInBuf[229]));
    OR3 i2_adj_56 (.O(n5239), .I0(n1_adj_281), .I1(state[0]), .I2(n2_adj_282));
    OR2 select_163_Select_163_i9 (.O(n9_adj_268), .I0(n2_adj_267), .I1(n1_adj_266));
    OR2 i3388 (.O(n6209), .I0(n6208), .I1(n6207));
    OR3 i1_adj_57 (.O(n5713), .I0(n1_adj_338), .I1(n2_adj_339), .I2(state[0]));
    AND2 select_163_Select_163_i2 (.O(n2_adj_267), .I0(state[6]), .I1(dataInBuf[155]));
    AND2 i3390 (.O(n6211), .I0(lcdRs_N_619), .I1(dataInBuf[230]));
    OR2 i3391 (.O(n6212), .I0(n6211), .I1(n6210));
    OR3 i2_adj_58 (.O(n5222), .I0(n1_adj_269), .I1(n2_adj_270), .I2(state[0]));
    OR3 i2_adj_59 (.O(n5242), .I0(n1_adj_260), .I1(state[0]), .I2(n2_adj_261));
    AND2 select_163_Select_162_i2 (.O(n2_adj_265), .I0(state[6]), .I1(dataInBuf[154]));
    AND2 i3393 (.O(n6214), .I0(lcdRs_N_619), .I1(dataInBuf[232]));
    AND2 i3018 (.O(n5839), .I0(lcdRs_N_619), .I1(dataInBuf[89]));
    OR2 i3394 (.O(n6215), .I0(n6214), .I1(n6213));
    OR3 i2_adj_60 (.O(n5244), .I0(n1_adj_195), .I1(state[0]), .I2(n2_adj_196));
    OR3 i1_adj_61 (.O(n5715), .I0(n1_adj_358), .I1(n2_adj_359), .I2(state[0]));
    AND2 select_163_Select_161_i2 (.O(n2_adj_263), .I0(state[6]), .I1(dataInBuf[153]));
    OR2 i3019 (.O(n5840), .I0(n5839), .I1(n5838));
    AND2 i3021 (.O(n5842), .I0(lcdRs_N_619), .I1(dataInBuf[90]));
    AND2 i3396 (.O(n6217), .I0(lcdRs_N_619), .I1(dataInBuf[233]));
    OR3 i2_adj_62 (.O(n5246), .I0(n1_adj_135), .I1(state[0]), .I2(n2_adj_136));
    OR2 i3397 (.O(n6218), .I0(n6217), .I1(n6216));
    AND2 i3399 (.O(n6220), .I0(lcdRs_N_619), .I1(dataInBuf[234]));
    OR3 i2_adj_63 (.O(n5248), .I0(n1_adj_91), .I1(state[0]), .I2(n2_adj_92));
    OR2 i3022 (.O(n5843), .I0(n5842), .I1(n5841));
    AND2 select_163_Select_160_i2 (.O(n2_adj_261), .I0(state[6]), .I1(dataInBuf[152]));
    OR2 i3400 (.O(n6221), .I0(n6220), .I1(n6219));
    AND2 i3024 (.O(n5845), .I0(lcdRs_N_619), .I1(dataInBuf[91]));
    AND2 i3402 (.O(n6223), .I0(lcdRs_N_619), .I1(dataInBuf[235]));
    OR2 i3403 (.O(n6224), .I0(n6223), .I1(n6222));
    OR3 i1_adj_64 (.O(lcdRs_N_618), .I0(dispCount[5]), .I1(n3800), .I2(n5));
    OR2 i3025 (.O(n5846), .I0(n5845), .I1(n5844));
    AND2 i3405 (.O(n6226), .I0(lcdRs_N_619), .I1(dataInBuf[236]));
    AND2 i3027 (.O(n5848), .I0(lcdRs_N_619), .I1(dataInBuf[92]));
    OR2 i3406 (.O(n6227), .I0(n6226), .I1(n6225));
    OR2 select_163_Select_158_i9 (.O(n9_adj_259), .I0(n2_adj_258), .I1(n1_adj_257));
    OR3 i1_adj_65 (.O(n5717), .I0(n1_adj_393), .I1(n2_adj_394), .I2(state[0]));
    OR2 i3028 (.O(n5849), .I0(n5848), .I1(n5847));
    AND2 i3408 (.O(n6229), .I0(lcdRs_N_619), .I1(dataInBuf[237]));
    AND2 i3030 (.O(n5851), .I0(lcdRs_N_619), .I1(dataInBuf[93]));
    AND2 select_163_Select_158_i2 (.O(n2_adj_258), .I0(state[6]), .I1(dataInBuf[150]));
    OR2 i3409 (.O(n6230), .I0(n6229), .I1(n6228));
    AND2 i3411 (.O(n6232), .I0(lcdRs_N_619), .I1(dataInBuf[238]));
    OR2 i3031 (.O(n5852), .I0(n5851), .I1(n5850));
    AND2 i3033 (.O(n5854), .I0(lcdRs_N_619), .I1(dataInBuf[94]));
    XOR2 i2912 (.O(n5733), .I0(dispCount[4]), .I1(dispCount[5]));
    OR2 i3412 (.O(n6233), .I0(n6232), .I1(n6231));
    OR2 i3034 (.O(n5855), .I0(n5854), .I1(n5853));
    AND2 select_163_Select_157_i2 (.O(n2_adj_256), .I0(state[6]), .I1(dataInBuf[149]));
    AND2 i3414 (.O(n6235), .I0(lcdRs_N_619), .I1(dataInBuf[240]));
    AND2 i3014 (.O(n5835), .I0(lcdRs_N_618), .I1(dataInBuf[80]));
    AND2 i3011 (.O(n5832), .I0(lcdRs_N_618), .I1(dataInBuf[78]));
    AND3 i2915 (.O(n3805), .I0(reset_c), .I1(n3649), .I2(n5735));
    AND2 i3008 (.O(n5829), .I0(lcdRs_N_618), .I1(dataInBuf[77]));
    OR2 i3415 (.O(n6236), .I0(n6235), .I1(n6234));
    OR2 i3424 (.O(n6245), .I0(n6244), .I1(n6243));
    OR2 i2923 (.O(n5744), .I0(n5743), .I1(n5742));
    AND2 i3005 (.O(n5826), .I0(lcdRs_N_618), .I1(dataInBuf[74]));
    OR2 select_163_Select_156_i9 (.O(n9_adj_254), .I0(n2_adj_253), .I1(n1_adj_252));
    AND2 i3002 (.O(n5823), .I0(lcdRs_N_618), .I1(dataInBuf[73]));
    OR2 select_163_Select_154_i9 (.O(n9_adj_248), .I0(n2_adj_247), .I1(n1_adj_246));
    OR2 i3037 (.O(n5858), .I0(n5857), .I1(n5856));
    AND2 i3426 (.O(n6247), .I0(lcdRs_N_619), .I1(dataInBuf[244]));
    OR2 i3427 (.O(n6248), .I0(n6247), .I1(n6246));
    AND2 i3039 (.O(n5860), .I0(lcdRs_N_619), .I1(dataInBuf[97]));
    AND2 select_163_Select_154_i2 (.O(n2_adj_247), .I0(state[6]), .I1(dataInBuf[146]));
    AND2 i3429 (.O(n6250), .I0(lcdRs_N_619), .I1(dataInBuf[245]));
    OR2 i3430 (.O(n6251), .I0(n6250), .I1(n6249));
    OR2 select_163_Select_153_i9 (.O(n9_adj_245), .I0(n2_adj_244), .I1(n1_adj_243));
    OR2 i3040 (.O(n5861), .I0(n5860), .I1(n5859));
    AND2 i3432 (.O(n6253), .I0(lcdRs_N_619), .I1(dataInBuf[246]));
    AND2 i3042 (.O(n5863), .I0(lcdRs_N_619), .I1(dataInBuf[98]));
    AND2 select_163_Select_153_i2 (.O(n2_adj_244), .I0(state[6]), .I1(dataInBuf[145]));
    OR2 i3433 (.O(n6254), .I0(n6253), .I1(n6252));
    AND2 i2999 (.O(n5820), .I0(lcdRs_N_618), .I1(dataInBuf[72]));
    AND2 i3435 (.O(n6256), .I0(lcdRs_N_619), .I1(dataInBuf[248]));
    OR2 i3043 (.O(n5864), .I0(n5863), .I1(n5862));
    OR2 select_163_Select_152_i9 (.O(n9_adj_242), .I0(n2_adj_241), .I1(n1_adj_240));
    OR2 i3436 (.O(n6257), .I0(n6256), .I1(n6255));
    AND2 i1_adj_66 (.O(n5719), .I0(n5718), .I1(state[1]));
    AND2 i3045 (.O(n5866), .I0(lcdRs_N_619), .I1(dataInBuf[99]));
    AND2 i3438 (.O(n6259), .I0(lcdRs_N_619), .I1(dataInBuf[249]));
    AND2 select_163_Select_152_i2 (.O(n2_adj_241), .I0(state[6]), .I1(dataInBuf[144]));
    OR2 i3439 (.O(n6260), .I0(n6259), .I1(n6258));
    AND2 i3441 (.O(n6262), .I0(lcdRs_N_619), .I1(dataInBuf[250]));
    AND2 i2996 (.O(n5817), .I0(lcdRs_N_618), .I1(dataInBuf[70]));
    OR2 i3442 (.O(n6263), .I0(n6262), .I1(n6261));
    OR3 i1_adj_67 (.O(n5669), .I0(n1_adj_93), .I1(n2_adj_94), .I2(state[0]));
    OR2 i3046 (.O(n5867), .I0(n5866), .I1(n5865));
    AND2 i3444 (.O(n6265), .I0(lcdRs_N_619), .I1(dataInBuf[251]));
    AND2 i3048 (.O(n5869), .I0(lcdRs_N_619), .I1(dataInBuf[100]));
    OR2 i3445 (.O(n6266), .I0(n6265), .I1(n6264));
    AND2 i3447 (.O(n6268), .I0(lcdRs_N_619), .I1(dataInBuf[252]));
    OR2 i3049 (.O(n5870), .I0(n5869), .I1(n5868));
    OR2 select_163_Select_150_i9 (.O(n9_adj_239), .I0(n2_adj_238), .I1(n1_adj_237));
    OR2 i3448 (.O(n6269), .I0(n6268), .I1(n6267));
    AND2 i3450 (.O(n6271), .I0(lcdRs_N_619), .I1(dataInBuf[253]));
    AND2 select_163_Select_150_i2 (.O(n2_adj_238), .I0(state[6]), .I1(dataInBuf[142]));
    AND2 i3051 (.O(n5872), .I0(lcdRs_N_619), .I1(dataInBuf[101]));
    OR2 i3451 (.O(n6272), .I0(n6271), .I1(n6270));
    AND2 i1_adj_68 (.O(n5720), .I0(lcdRs_N_619), .I1(state[7]));
    AND2 i3453 (.O(n6274), .I0(lcdRs_N_619), .I1(dataInBuf[254]));
    OR3 i1_adj_69 (.O(n1845), .I0(n1_adj_10), .I1(n3800), .I2(dispCount[4]));
    OR2 i3454 (.O(n6275), .I0(n6274), .I1(n6273));
    OR2 i3052 (.O(n5873), .I0(n5872), .I1(n5871));
    AND2 i3456 (.O(n6277), .I0(n2185), .I1(dataInBuf[250]));
    OR2 i3457 (.O(n6278), .I0(n6277), .I1(n6276));
    AND2 select_163_Select_149_i2 (.O(n2_adj_236), .I0(state[6]), .I1(dataInBuf[141]));
    AND2 i3054 (.O(n5875), .I0(lcdRs_N_619), .I1(dataInBuf[102]));
    AND2 i3459 (.O(n6280), .I0(n2185), .I1(dataInBuf[249]));
    OR2 select_163_Select_148_i9 (.O(n9_adj_234), .I0(n2_adj_233), .I1(n1_adj_232));
    OR2 i3055 (.O(n5876), .I0(n5875), .I1(n5874));
    AND2 i1_adj_70 (.O(n5721), .I0(n5720), .I1(dataInBuf[34]));
    OR2 i3460 (.O(n6281), .I0(n6280), .I1(n6279));
    AND2 i3462 (.O(n6283), .I0(n2185), .I1(dataInBuf[248]));
    AND2 select_163_Select_148_i2 (.O(n2_adj_233), .I0(state[6]), .I1(dataInBuf[140]));
    OR2 i3463 (.O(n6284), .I0(n6283), .I1(n6282));
    AND2 i2276 (.O(n5099), .I0(n5092), .I1(cnt[7]));
    OR2 select_163_Select_147_i9 (.O(n9_adj_231), .I0(n2_adj_230), .I1(n1_adj_229));
    OR3 i1_adj_71 (.O(n5671), .I0(n1_adj_155), .I1(n2_adj_156), .I2(state[0]));
    AND2 i1_adj_72 (.O(n3644), .I0(n5720), .I1(n1845));
    AND2 i3057 (.O(n5878), .I0(lcdRs_N_619), .I1(dataInBuf[104]));
    AND2 i3465 (.O(n6286), .I0(n6285), .I1(n44));
    AND2 select_163_Select_147_i2 (.O(n2_adj_230), .I0(state[6]), .I1(dataInBuf[139]));
    AND3 i3466 (.O(n6287), .I0(n2185), .I1(n60), .I2(dataInBuf[253]));
    OR2 i3467 (.O(n6288), .I0(n6287), .I1(n6286));
    OR2 i3058 (.O(n5879), .I0(n5878), .I1(n5877));
    OR2 select_163_Select_146_i9 (.O(n9_adj_228), .I0(n2_adj_227), .I1(n1_adj_226));
    AND3 i3469 (.O(n6290), .I0(n2185), .I1(n60), .I2(dataInBuf[252]));
    AND2 i3060 (.O(n5881), .I0(lcdRs_N_619), .I1(dataInBuf[105]));
    OR2 i3470 (.O(n6291), .I0(n6290), .I1(n6289));
    AND2 select_163_Select_146_i2 (.O(n2_adj_227), .I0(state[6]), .I1(dataInBuf[138]));
    AND3 i3472 (.O(n6293), .I0(n2185), .I1(n60), .I2(dataInBuf[251]));
    OR2 i3061 (.O(n5882), .I0(n5881), .I1(n5880));
    OR2 select_163_Select_145_i9 (.O(n9_adj_225), .I0(n2_adj_224), .I1(n1_adj_223));
    OR2 i3473 (.O(n6294), .I0(n6293), .I1(n6292));
    XOR2 i2259 (.O(n100), .I0(n5078), .I1(cnt[5]));
    AND2 i3063 (.O(n5884), .I0(lcdRs_N_619), .I1(dataInBuf[106]));
    AND2 select_163_Select_145_i2 (.O(n2_adj_224), .I0(state[6]), .I1(dataInBuf[137]));
    OR2 select_163_Select_144_i9 (.O(n9_adj_222), .I0(n2_adj_221), .I1(n1_adj_220));
    OR2 i3064 (.O(n5885), .I0(n5884), .I1(n5883));
    OR3 i1_adj_73 (.O(n5673), .I0(n2_adj_396), .I1(n1_adj_395), .I2(state[0]));
    AND2 select_163_Select_144_i2 (.O(n2_adj_221), .I0(state[6]), .I1(dataInBuf[136]));
    AND2 i3066 (.O(n5887), .I0(lcdRs_N_619), .I1(dataInBuf[107]));
    OR2 i3067 (.O(n5888), .I0(n5887), .I1(n5886));
    AND2 i3069 (.O(n5890), .I0(lcdRs_N_619), .I1(dataInBuf[108]));
    OR2 i3070 (.O(n5891), .I0(n5890), .I1(n5889));
    OR2 select_163_Select_142_i9 (.O(n9_adj_219), .I0(n2_adj_218), .I1(n1_adj_217));
    AND2 i3072 (.O(n5893), .I0(lcdRs_N_619), .I1(dataInBuf[109]));
    OR2 i3073 (.O(n5894), .I0(n5893), .I1(n5892));
    AND2 select_163_Select_142_i2 (.O(n2_adj_218), .I0(state[6]), .I1(dataInBuf[134]));
    AND2 i3075 (.O(n5896), .I0(lcdRs_N_619), .I1(dataInBuf[110]));
    OR2 i3076 (.O(n5897), .I0(n5896), .I1(n5895));
    AND2 select_163_Select_141_i2 (.O(n2_adj_216), .I0(state[6]), .I1(dataInBuf[133]));
    OR2 select_163_Select_140_i9 (.O(n9_adj_214), .I0(n2_adj_213), .I1(n1_adj_212));
    AND2 i2993 (.O(n5814), .I0(lcdRs_N_618), .I1(dataInBuf[69]));
    AND2 i1_adj_74 (.O(n5723), .I0(n5720), .I1(dataInBuf[83]));
    AND2 i3078 (.O(n5899), .I0(lcdRs_N_619), .I1(dataInBuf[112]));
    AND2 select_163_Select_140_i2 (.O(n2_adj_213), .I0(state[6]), .I1(dataInBuf[132]));
    OR2 select_163_Select_139_i9 (.O(n9_adj_211), .I0(n2_adj_210), .I1(n1_adj_209));
    OR2 i3079 (.O(n5900), .I0(n5899), .I1(n5898));
    AND2 i3081 (.O(n5902), .I0(lcdRs_N_619), .I1(dataInBuf[113]));
    AND2 select_163_Select_139_i2 (.O(n2_adj_210), .I0(state[6]), .I1(dataInBuf[131]));
    OR2 i3082 (.O(n5903), .I0(n5902), .I1(n5901));
    OR2 select_163_Select_138_i9 (.O(n9_adj_208), .I0(n2_adj_207), .I1(n1_adj_206));
    AND2 i3084 (.O(n5905), .I0(lcdRs_N_619), .I1(dataInBuf[114]));
    AND2 i2990 (.O(n5811), .I0(lcdRs_N_618), .I1(dataInBuf[66]));
    AND2 i1_adj_75 (.O(n5724), .I0(n5720), .I1(dataInBuf[5]));
    AND2 select_163_Select_138_i2 (.O(n2_adj_207), .I0(state[6]), .I1(dataInBuf[130]));
    OR2 select_163_Select_137_i9 (.O(n9_adj_205), .I0(n2_adj_204), .I1(n1_adj_203));
    OR3 i1_adj_76 (.O(n5675), .I0(n2_adj_377), .I1(n1_adj_376), .I2(state[0]));
    XOR2 i2266 (.O(n99), .I0(n5085), .I1(cnt[6]));
    OR2 i3085 (.O(n5906), .I0(n5905), .I1(n5904));
    AND2 select_163_Select_137_i2 (.O(n2_adj_204), .I0(state[6]), .I1(dataInBuf[129]));
    AND2 i3087 (.O(n5908), .I0(lcdRs_N_619), .I1(dataInBuf[115]));
    OR2 select_163_Select_136_i9 (.O(n9_adj_202), .I0(n2_adj_201), .I1(n1_adj_200));
    OR2 i3088 (.O(n5909), .I0(n5908), .I1(n5907));
    AND2 i1_adj_77 (.O(n5725), .I0(n5720), .I1(dataInBuf[38]));
    AND2 select_163_Select_136_i2 (.O(n2_adj_201), .I0(state[6]), .I1(dataInBuf[128]));
    AND2 i1_adj_78 (.O(n5726), .I0(n5720), .I1(dataInBuf[48]));
    XOR2 i2273 (.O(n98), .I0(n5092), .I1(cnt[7]));
    AND2 i3090 (.O(n5911), .I0(lcdRs_N_619), .I1(dataInBuf[116]));
    XOR2 i2280 (.O(n97), .I0(n5099), .I1(cnt[8]));
    OR2 i3091 (.O(n5912), .I0(n5911), .I1(n5910));
    OR2 select_163_Select_134_i9 (.O(n9_adj_199), .I0(n2_adj_198), .I1(n1_adj_197));
    AND2 i3093 (.O(n5914), .I0(lcdRs_N_619), .I1(dataInBuf[117]));
    OR2 i3094 (.O(n5915), .I0(n5914), .I1(n5913));
    AND2 select_163_Select_134_i2 (.O(n2_adj_198), .I0(state[6]), .I1(dataInBuf[126]));
    AND2 i3096 (.O(n5917), .I0(lcdRs_N_619), .I1(dataInBuf[118]));
    AND2 select_163_Select_133_i2 (.O(n2_adj_196), .I0(state[6]), .I1(dataInBuf[125]));
    OR2 i3097 (.O(n5918), .I0(n5917), .I1(n5916));
    AND2 i3099 (.O(n5920), .I0(lcdRs_N_619), .I1(dataInBuf[120]));
    OR2 select_163_Select_132_i9 (.O(n9_adj_194), .I0(n2_adj_193), .I1(n1_adj_192));
    AND2 i1_adj_79 (.O(n5727), .I0(n5720), .I1(dataInBuf[33]));
    AND2 select_163_Select_132_i2 (.O(n2_adj_193), .I0(state[6]), .I1(dataInBuf[124]));
    OR2 i3100 (.O(n5921), .I0(n5920), .I1(n5919));
    OR2 select_163_Select_131_i9 (.O(n9_adj_191), .I0(n2_adj_190), .I1(n1_adj_189));
    OR3 i1_adj_80 (.O(n5677), .I0(n2_adj_357), .I1(n1_adj_356), .I2(state[0]));
    AND2 i3102 (.O(n5923), .I0(lcdRs_N_619), .I1(dataInBuf[121]));
    XOR2 i2287 (.O(n96), .I0(n5106), .I1(cnt[9]));
    AND2 select_163_Select_131_i2 (.O(n2_adj_190), .I0(state[6]), .I1(dataInBuf[123]));
    AND2 i1_adj_81 (.O(n5728), .I0(n5720), .I1(dataInBuf[84]));
    OR2 select_163_Select_130_i9 (.O(n9_adj_188), .I0(n2_adj_187), .I1(n1_adj_186));
    OR2 i3103 (.O(n5924), .I0(n5923), .I1(n5922));
    AND2 select_163_Select_130_i2 (.O(n2_adj_187), .I0(state[6]), .I1(dataInBuf[122]));
    OR2 select_163_Select_129_i9 (.O(n9_adj_185), .I0(n2_adj_184), .I1(n1_adj_183));
    AND2 i3105 (.O(n5926), .I0(lcdRs_N_619), .I1(dataInBuf[122]));
    AND2 select_163_Select_129_i2 (.O(n2_adj_184), .I0(state[6]), .I1(dataInBuf[121]));
    OR2 select_163_Select_128_i9 (.O(n9_adj_182), .I0(n2_adj_181), .I1(n1_adj_180));
    OR2 i3106 (.O(n5927), .I0(n5926), .I1(n5925));
    AND2 i3108 (.O(n5929), .I0(lcdRs_N_619), .I1(dataInBuf[123]));
    AND2 select_163_Select_128_i2 (.O(n2_adj_181), .I0(state[6]), .I1(dataInBuf[120]));
    OR3 i1_adj_82 (.O(n5679), .I0(n2_adj_331), .I1(n1_adj_330), .I2(state[0]));
    OR2 i3109 (.O(n5930), .I0(n5929), .I1(n5928));
    XOR2 i2294 (.O(n95), .I0(n5113), .I1(cnt[10]));
    OR2 select_163_Select_126_i9 (.O(n9_adj_179), .I0(n2_adj_178), .I1(n1_adj_177));
    AND2 i3111 (.O(n5932), .I0(lcdRs_N_619), .I1(dataInBuf[124]));
    AND2 select_163_Select_126_i2 (.O(n2_adj_178), .I0(state[6]), .I1(dataInBuf[118]));
    OR2 i3112 (.O(n5933), .I0(n5932), .I1(n5931));
    AND2 i3114 (.O(n5935), .I0(lcdRs_N_619), .I1(dataInBuf[125]));
    OR2 i3115 (.O(n5936), .I0(n5935), .I1(n5934));
    AND2 select_163_Select_125_i2 (.O(n2_adj_176), .I0(state[6]), .I1(dataInBuf[117]));
    AND2 i2987 (.O(n5808), .I0(lcdRs_N_618), .I1(dataInBuf[65]));
    AND2 i3117 (.O(n5938), .I0(lcdRs_N_619), .I1(dataInBuf[126]));
    AND2 i3189 (.O(n6010), .I0(lcdRs_N_619), .I1(dataInBuf[154]));
    AND2 i2984 (.O(n5805), .I0(lcdRs_N_618), .I1(dataInBuf[64]));
    AND2 i2981 (.O(n5802), .I0(lcdRs_N_618), .I1(dataInBuf[62]));
    AND2 i2978 (.O(n5799), .I0(lcdRs_N_618), .I1(dataInBuf[61]));
    AND2 i2975 (.O(n5796), .I0(lcdRs_N_618), .I1(dataInBuf[58]));
    AND2 i2972 (.O(n5793), .I0(lcdRs_N_618), .I1(dataInBuf[57]));
    AND2 i2969 (.O(n5790), .I0(lcdRs_N_618), .I1(dataInBuf[56]));
    AND2 i2966 (.O(n5787), .I0(lcdRs_N_618), .I1(dataInBuf[54]));
    AND2 i2963 (.O(n5784), .I0(lcdRs_N_618), .I1(dataInBuf[53]));
    AND2 i2960 (.O(n5781), .I0(lcdRs_N_618), .I1(dataInBuf[50]));
    AND2 i2957 (.O(n5778), .I0(lcdRs_N_618), .I1(dataInBuf[49]));
    AND2 i2954 (.O(n5775), .I0(lcdRs_N_618), .I1(dataInBuf[48]));
    AND2 i2951 (.O(n5772), .I0(lcdRs_N_618), .I1(dataInBuf[46]));
    AND2 i2318 (.O(n5141), .I0(n5134), .I1(cnt[13]));
    INV i2914 (.O(n5735), .I0(n2212));
    INV i2229 (.O(n105), .I0(cnt[0]));
    AND2 i1_adj_83 (.O(n21), .I0(cnt[18]), .I1(cnt[7]));
    OR3 i1_adj_84 (.O(n5689), .I0(n2_adj_265), .I1(n1_adj_264), .I2(state[0]));
    AND2 i2948 (.O(n5769), .I0(lcdRs_N_618), .I1(dataInBuf[45]));
    INV i3464 (.O(n6285), .I0(n60));
    INV i264 (.O(n14_adj_6), .I0(state[3]));
    INV i1598 (.O(n3729), .I0(n3800));
    AND2 i2945 (.O(n5766), .I0(lcdRs_N_618), .I1(dataInBuf[42]));
    OR3 i2_adj_85 (.O(n5216), .I0(n1_adj_328), .I1(n2_adj_329), .I2(state[0]));
    INV i2908 (.O(n5718), .I0(n5729));
    INV i979 (.O(n3806), .I0(n2212));
    VCC i2911 (.X(pwr));
    AND2 i2942 (.O(n5763), .I0(lcdRs_N_618), .I1(dataInBuf[41]));
    AND2 i2939 (.O(n5760), .I0(lcdRs_N_618), .I1(dataInBuf[38]));
    AND2 i6 (.O(n26), .I0(cnt[1]), .I1(cnt[17]));
    AND2 i7 (.O(n27), .I0(cnt[10]), .I1(cnt[5]));
    AND2 i8 (.O(n28), .I0(cnt[4]), .I1(cnt[19]));
    AND2 i2936 (.O(n5757), .I0(lcdRs_N_618), .I1(dataInBuf[37]));
    AND2 i2933 (.O(n5754), .I0(lcdRs_N_618), .I1(dataInBuf[34]));
    AND2 i9 (.O(n29), .I0(cnt[15]), .I1(cnt[12]));
    INV i1551 (.O(n4376), .I0(n3012));
    AND2 i10 (.O(n30), .I0(cnt[11]), .I1(cnt[2]));
    AND2 i2325 (.O(n5148), .I0(n5141), .I1(cnt[14]));
    OR3 i2_adj_86 (.O(n5214), .I0(n1_adj_348), .I1(n2_adj_349), .I2(state[0]));
    INV i1549 (.O(n4374), .I0(n2185));
    AND2 i11 (.O(n31), .I0(n22), .I1(n21));
    AND2 i12 (.O(n32), .I0(n24), .I1(n23));
    AND2 i2930 (.O(n5751), .I0(lcdRs_N_618), .I1(dataInBuf[33]));
    OR3 i2_adj_87 (.O(n5212), .I0(n1_adj_374), .I1(n2_adj_375), .I2(state[0]));
    INV equal_76_i12 (.O(lcdRs_N_619), .I0(lcdRs_N_618));
    INV i2913 (.O(n5734), .I0(n5733));
    INV i1_adj_88 (.O(n1_adj_10), .I0(dispCount[5]));
    OR2 i3190 (.O(n6011), .I0(n6010), .I1(n6009));
    AND2 i2927 (.O(n5748), .I0(lcdRs_N_618), .I1(dataInBuf[29]));
    INV equal_75_i12 (.O(lcdRs_N_620), .I0(n1845));
    INV i15 (.O(n3006), .I0(n14));
    INV i6_adj_89 (.O(dispCount_5__N_347[0]), .I0(dispCount[0]));
    AND2 i3192 (.O(n6013), .I0(lcdRs_N_619), .I1(dataInBuf[155]));
    AND2 i2924 (.O(n5745), .I0(lcdRs_N_618), .I1(dataInBuf[21]));
    INV i1_adj_90 (.O(n1), .I0(state[7]));
    AND2 i14 (.O(n34), .I0(n28), .I1(n27));
    AND2 i15_adj_91 (.O(n35), .I0(n30), .I1(n29));
    OR2 i3193 (.O(n6014), .I0(n6013), .I1(n6012));
    AND2 i3195 (.O(n6016), .I0(lcdRs_N_619), .I1(dataInBuf[156]));
    AND2 i2_adj_92 (.O(n22), .I0(cnt[3]), .I1(cnt[16]));
    AND2 i16 (.O(n36), .I0(n32), .I1(n31));
    AND2 i3_adj_93 (.O(n23), .I0(cnt[0]), .I1(cnt[6]));
    AND2 i2921 (.O(n5742), .I0(lcdRs_N_618), .I1(dataInBuf[13]));
    INV i1594 (.O(n3100), .I0(n5258));
    INV i229 (.O(n5), .I0(dispCount[4]));
    DFFR state_FSM_i6 (.Q(state[1]), .D(state[0]), .CLK(ledEN_c), .R(reset_c));   // lcd1602.v(63[13] 138[20])
    DFFR state_FSM_i5 (.Q(state[2]), .D(state[1]), .CLK(ledEN_c), .R(reset_c));   // lcd1602.v(63[13] 138[20])
    DFFR state_FSM_i4 (.Q(state[3]), .D(state[2]), .CLK(ledEN_c), .R(reset_c));   // lcd1602.v(63[13] 138[20])
    DFFR state_FSM_i3 (.Q(state[4]), .D(state[3]), .CLK(ledEN_c), .R(reset_c));   // lcd1602.v(63[13] 138[20])
    DFFR state_FSM_i2 (.Q(state[6]), .D(n3644), .CLK(ledEN_c), .R(reset_c));   // lcd1602.v(63[13] 138[20])
    DFFCR dispCount_i0_i5 (.Q(dispCount[5]), .D(n2164), .CLK(ledEN_c), 
          .CE(n3804), .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR dispCount_i0_i4 (.Q(dispCount[4]), .D(n2163), .CLK(ledEN_c), 
          .CE(n3804), .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR dispCount_i0_i3 (.Q(dispCount[3]), .D(n2162), .CLK(ledEN_c), 
          .CE(n3804), .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR dispCount_i0_i2 (.Q(dispCount[2]), .D(n2161), .CLK(ledEN_c), 
          .CE(n3804), .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR dispCount_i0_i1 (.Q(dispCount[1]), .D(n2160), .CLK(ledEN_c), 
          .CE(n3804), .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR lcdD_i0_i8 (.Q(lcdD_c_7), .D(n3638), .CLK(ledEN_c), .CE(n3806), 
          .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR lcdD_i0_i7 (.Q(lcdD_c_6), .D(n2199), .CLK(ledEN_c), .CE(n3806), 
          .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR lcdD_i0_i6 (.Q(lcdD_c_5), .D(n6288), .CLK(ledEN_c), .CE(n3806), 
          .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR lcdD_i0_i5 (.Q(lcdD_c_4), .D(n6291), .CLK(ledEN_c), .CE(n3806), 
          .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR lcdD_i0_i4 (.Q(lcdD_c_3), .D(n6294), .CLK(ledEN_c), .CE(n3806), 
          .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR lcdD_i0_i3 (.Q(lcdD_c_2), .D(n6278), .CLK(ledEN_c), .CE(n3806), 
          .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCR lcdD_i0_i2 (.Q(lcdD_c_1), .D(n6281), .CLK(ledEN_c), .CE(n3806), 
          .R(reset_c));   // lcd1602.v(62[14] 139[12])
    DFFCS lcdD_i0_i1 (.Q(lcdD_c_0), .D(n6284), .CLK(ledEN_c), .CE(n3806), 
          .S(reset_c));   // lcd1602.v(62[14] 139[12])
    OBUF lcdD_pad_6 (.O(lcdD[6]), .I0(lcdD_c_6));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    IBUF clk_50m_pad (.O(clk_50m_c), .I0(clk_50m));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(186[8:12])
    OBUF ledEN_pad (.O(ledEN), .I0(ledEN_c));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF lcdRw_pad (.O(lcdRw), .I0(lcdRw_c));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF lcdRs_pad (.O(lcdRs), .I0(lcdRs_c));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF lcdD_pad_0 (.O(lcdD[0]), .I0(lcdD_c_0));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF lcdD_pad_1 (.O(lcdD[1]), .I0(lcdD_c_1));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF lcdD_pad_2 (.O(lcdD[2]), .I0(lcdD_c_2));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF lcdD_pad_3 (.O(lcdD[3]), .I0(lcdD_c_3));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF lcdD_pad_4 (.O(lcdD[4]), .I0(lcdD_c_4));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    OBUF lcdD_pad_5 (.O(lcdD[5]), .I0(lcdD_c_5));   // D:/ispLEVER_Classic2_1/lse/userware/NT/SYNTHESIS_HEADERS/mach.v(270[8:12])
    AND2 i4 (.O(n24), .I0(cnt[14]), .I1(cnt[9]));
    
endmodule
//
// Verilog Description of module GND
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR2
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND2
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR3
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND3
// module not written out since it is a black-box. 
//

//
// Verilog Description of module INV
// module not written out since it is a black-box. 
//

//
// Verilog Description of module XOR2
// module not written out since it is a black-box. 
//

//
// Verilog Description of module OR4
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND6
// module not written out since it is a black-box. 
//

//
// Verilog Description of module AND4
// module not written out since it is a black-box. 
//

//
// Verilog Description of module VCC
// module not written out since it is a black-box. 
//

